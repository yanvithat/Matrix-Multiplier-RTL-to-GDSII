module matrix_mult3 (clk,
    input_a_serial,
    input_b_serial,
    rst,
    output_c_serial);
 input clk;
 input input_a_serial;
 input input_b_serial;
 input rst;
 output [31:0] output_c_serial;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire \input_a[0][0] ;
 wire \input_a[10][0] ;
 wire \input_a[11][0] ;
 wire \input_a[12][0] ;
 wire \input_a[13][0] ;
 wire \input_a[14][0] ;
 wire \input_a[15] ;
 wire \input_a[1][0] ;
 wire \input_a[2][0] ;
 wire \input_a[3][0] ;
 wire \input_a[4][0] ;
 wire \input_a[5][0] ;
 wire \input_a[6][0] ;
 wire \input_a[7][0] ;
 wire \input_a[8][0] ;
 wire \input_a[9][0] ;
 wire \input_b[15][0] ;
 wire \output_c[0][0] ;
 wire \output_c[0][10] ;
 wire \output_c[0][11] ;
 wire \output_c[0][12] ;
 wire \output_c[0][13] ;
 wire \output_c[0][14] ;
 wire \output_c[0][15] ;
 wire \output_c[0][16] ;
 wire \output_c[0][17] ;
 wire \output_c[0][18] ;
 wire \output_c[0][19] ;
 wire \output_c[0][1] ;
 wire \output_c[0][20] ;
 wire \output_c[0][21] ;
 wire \output_c[0][22] ;
 wire \output_c[0][23] ;
 wire \output_c[0][24] ;
 wire \output_c[0][25] ;
 wire \output_c[0][26] ;
 wire \output_c[0][27] ;
 wire \output_c[0][28] ;
 wire \output_c[0][29] ;
 wire \output_c[0][2] ;
 wire \output_c[0][30] ;
 wire \output_c[0][31] ;
 wire \output_c[0][3] ;
 wire \output_c[0][4] ;
 wire \output_c[0][5] ;
 wire \output_c[0][6] ;
 wire \output_c[0][7] ;
 wire \output_c[0][8] ;
 wire \output_c[0][9] ;
 wire \output_c[10][0] ;
 wire \output_c[10][10] ;
 wire \output_c[10][11] ;
 wire \output_c[10][12] ;
 wire \output_c[10][13] ;
 wire \output_c[10][14] ;
 wire \output_c[10][15] ;
 wire \output_c[10][16] ;
 wire \output_c[10][17] ;
 wire \output_c[10][18] ;
 wire \output_c[10][19] ;
 wire \output_c[10][1] ;
 wire \output_c[10][20] ;
 wire \output_c[10][21] ;
 wire \output_c[10][22] ;
 wire \output_c[10][23] ;
 wire \output_c[10][24] ;
 wire \output_c[10][25] ;
 wire \output_c[10][26] ;
 wire \output_c[10][27] ;
 wire \output_c[10][28] ;
 wire \output_c[10][29] ;
 wire \output_c[10][2] ;
 wire \output_c[10][30] ;
 wire \output_c[10][31] ;
 wire \output_c[10][3] ;
 wire \output_c[10][4] ;
 wire \output_c[10][5] ;
 wire \output_c[10][6] ;
 wire \output_c[10][7] ;
 wire \output_c[10][8] ;
 wire \output_c[10][9] ;
 wire \output_c[11][0] ;
 wire \output_c[11][10] ;
 wire \output_c[11][11] ;
 wire \output_c[11][12] ;
 wire \output_c[11][13] ;
 wire \output_c[11][14] ;
 wire \output_c[11][15] ;
 wire \output_c[11][16] ;
 wire \output_c[11][17] ;
 wire \output_c[11][18] ;
 wire \output_c[11][19] ;
 wire \output_c[11][1] ;
 wire \output_c[11][20] ;
 wire \output_c[11][21] ;
 wire \output_c[11][22] ;
 wire \output_c[11][23] ;
 wire \output_c[11][24] ;
 wire \output_c[11][25] ;
 wire \output_c[11][26] ;
 wire \output_c[11][27] ;
 wire \output_c[11][28] ;
 wire \output_c[11][29] ;
 wire \output_c[11][2] ;
 wire \output_c[11][30] ;
 wire \output_c[11][31] ;
 wire \output_c[11][3] ;
 wire \output_c[11][4] ;
 wire \output_c[11][5] ;
 wire \output_c[11][6] ;
 wire \output_c[11][7] ;
 wire \output_c[11][8] ;
 wire \output_c[11][9] ;
 wire \output_c[12][0] ;
 wire \output_c[12][10] ;
 wire \output_c[12][11] ;
 wire \output_c[12][12] ;
 wire \output_c[12][13] ;
 wire \output_c[12][14] ;
 wire \output_c[12][15] ;
 wire \output_c[12][16] ;
 wire \output_c[12][17] ;
 wire \output_c[12][18] ;
 wire \output_c[12][19] ;
 wire \output_c[12][1] ;
 wire \output_c[12][20] ;
 wire \output_c[12][21] ;
 wire \output_c[12][22] ;
 wire \output_c[12][23] ;
 wire \output_c[12][24] ;
 wire \output_c[12][25] ;
 wire \output_c[12][26] ;
 wire \output_c[12][27] ;
 wire \output_c[12][28] ;
 wire \output_c[12][29] ;
 wire \output_c[12][2] ;
 wire \output_c[12][30] ;
 wire \output_c[12][31] ;
 wire \output_c[12][3] ;
 wire \output_c[12][4] ;
 wire \output_c[12][5] ;
 wire \output_c[12][6] ;
 wire \output_c[12][7] ;
 wire \output_c[12][8] ;
 wire \output_c[12][9] ;
 wire \output_c[13][0] ;
 wire \output_c[13][10] ;
 wire \output_c[13][11] ;
 wire \output_c[13][12] ;
 wire \output_c[13][13] ;
 wire \output_c[13][14] ;
 wire \output_c[13][15] ;
 wire \output_c[13][16] ;
 wire \output_c[13][17] ;
 wire \output_c[13][18] ;
 wire \output_c[13][19] ;
 wire \output_c[13][1] ;
 wire \output_c[13][20] ;
 wire \output_c[13][21] ;
 wire \output_c[13][22] ;
 wire \output_c[13][23] ;
 wire \output_c[13][24] ;
 wire \output_c[13][25] ;
 wire \output_c[13][26] ;
 wire \output_c[13][27] ;
 wire \output_c[13][28] ;
 wire \output_c[13][29] ;
 wire \output_c[13][2] ;
 wire \output_c[13][30] ;
 wire \output_c[13][31] ;
 wire \output_c[13][3] ;
 wire \output_c[13][4] ;
 wire \output_c[13][5] ;
 wire \output_c[13][6] ;
 wire \output_c[13][7] ;
 wire \output_c[13][8] ;
 wire \output_c[13][9] ;
 wire \output_c[14][0] ;
 wire \output_c[14][10] ;
 wire \output_c[14][11] ;
 wire \output_c[14][12] ;
 wire \output_c[14][13] ;
 wire \output_c[14][14] ;
 wire \output_c[14][15] ;
 wire \output_c[14][16] ;
 wire \output_c[14][17] ;
 wire \output_c[14][18] ;
 wire \output_c[14][19] ;
 wire \output_c[14][1] ;
 wire \output_c[14][20] ;
 wire \output_c[14][21] ;
 wire \output_c[14][22] ;
 wire \output_c[14][23] ;
 wire \output_c[14][24] ;
 wire \output_c[14][25] ;
 wire \output_c[14][26] ;
 wire \output_c[14][27] ;
 wire \output_c[14][28] ;
 wire \output_c[14][29] ;
 wire \output_c[14][2] ;
 wire \output_c[14][30] ;
 wire \output_c[14][31] ;
 wire \output_c[14][3] ;
 wire \output_c[14][4] ;
 wire \output_c[14][5] ;
 wire \output_c[14][6] ;
 wire \output_c[14][7] ;
 wire \output_c[14][8] ;
 wire \output_c[14][9] ;
 wire \output_c[15][0] ;
 wire \output_c[15][10] ;
 wire \output_c[15][11] ;
 wire \output_c[15][12] ;
 wire \output_c[15][13] ;
 wire \output_c[15][14] ;
 wire \output_c[15][15] ;
 wire \output_c[15][16] ;
 wire \output_c[15][17] ;
 wire \output_c[15][18] ;
 wire \output_c[15][19] ;
 wire \output_c[15][1] ;
 wire \output_c[15][20] ;
 wire \output_c[15][21] ;
 wire \output_c[15][22] ;
 wire \output_c[15][23] ;
 wire \output_c[15][24] ;
 wire \output_c[15][25] ;
 wire \output_c[15][26] ;
 wire \output_c[15][27] ;
 wire \output_c[15][28] ;
 wire \output_c[15][29] ;
 wire \output_c[15][2] ;
 wire \output_c[15][30] ;
 wire \output_c[15][31] ;
 wire \output_c[15][3] ;
 wire \output_c[15][4] ;
 wire \output_c[15][5] ;
 wire \output_c[15][6] ;
 wire \output_c[15][7] ;
 wire \output_c[15][8] ;
 wire \output_c[15][9] ;
 wire \output_c[1][0] ;
 wire \output_c[1][10] ;
 wire \output_c[1][11] ;
 wire \output_c[1][12] ;
 wire \output_c[1][13] ;
 wire \output_c[1][14] ;
 wire \output_c[1][15] ;
 wire \output_c[1][16] ;
 wire \output_c[1][17] ;
 wire \output_c[1][18] ;
 wire \output_c[1][19] ;
 wire \output_c[1][1] ;
 wire \output_c[1][20] ;
 wire \output_c[1][21] ;
 wire \output_c[1][22] ;
 wire \output_c[1][23] ;
 wire \output_c[1][24] ;
 wire \output_c[1][25] ;
 wire \output_c[1][26] ;
 wire \output_c[1][27] ;
 wire \output_c[1][28] ;
 wire \output_c[1][29] ;
 wire \output_c[1][2] ;
 wire \output_c[1][30] ;
 wire \output_c[1][31] ;
 wire \output_c[1][3] ;
 wire \output_c[1][4] ;
 wire \output_c[1][5] ;
 wire \output_c[1][6] ;
 wire \output_c[1][7] ;
 wire \output_c[1][8] ;
 wire \output_c[1][9] ;
 wire \output_c[2][0] ;
 wire \output_c[2][10] ;
 wire \output_c[2][11] ;
 wire \output_c[2][12] ;
 wire \output_c[2][13] ;
 wire \output_c[2][14] ;
 wire \output_c[2][15] ;
 wire \output_c[2][16] ;
 wire \output_c[2][17] ;
 wire \output_c[2][18] ;
 wire \output_c[2][19] ;
 wire \output_c[2][1] ;
 wire \output_c[2][20] ;
 wire \output_c[2][21] ;
 wire \output_c[2][22] ;
 wire \output_c[2][23] ;
 wire \output_c[2][24] ;
 wire \output_c[2][25] ;
 wire \output_c[2][26] ;
 wire \output_c[2][27] ;
 wire \output_c[2][28] ;
 wire \output_c[2][29] ;
 wire \output_c[2][2] ;
 wire \output_c[2][30] ;
 wire \output_c[2][31] ;
 wire \output_c[2][3] ;
 wire \output_c[2][4] ;
 wire \output_c[2][5] ;
 wire \output_c[2][6] ;
 wire \output_c[2][7] ;
 wire \output_c[2][8] ;
 wire \output_c[2][9] ;
 wire \output_c[3][0] ;
 wire \output_c[3][10] ;
 wire \output_c[3][11] ;
 wire \output_c[3][12] ;
 wire \output_c[3][13] ;
 wire \output_c[3][14] ;
 wire \output_c[3][15] ;
 wire \output_c[3][16] ;
 wire \output_c[3][17] ;
 wire \output_c[3][18] ;
 wire \output_c[3][19] ;
 wire \output_c[3][1] ;
 wire \output_c[3][20] ;
 wire \output_c[3][21] ;
 wire \output_c[3][22] ;
 wire \output_c[3][23] ;
 wire \output_c[3][24] ;
 wire \output_c[3][25] ;
 wire \output_c[3][26] ;
 wire \output_c[3][27] ;
 wire \output_c[3][28] ;
 wire \output_c[3][29] ;
 wire \output_c[3][2] ;
 wire \output_c[3][30] ;
 wire \output_c[3][31] ;
 wire \output_c[3][3] ;
 wire \output_c[3][4] ;
 wire \output_c[3][5] ;
 wire \output_c[3][6] ;
 wire \output_c[3][7] ;
 wire \output_c[3][8] ;
 wire \output_c[3][9] ;
 wire \output_c[4][0] ;
 wire \output_c[4][10] ;
 wire \output_c[4][11] ;
 wire \output_c[4][12] ;
 wire \output_c[4][13] ;
 wire \output_c[4][14] ;
 wire \output_c[4][15] ;
 wire \output_c[4][16] ;
 wire \output_c[4][17] ;
 wire \output_c[4][18] ;
 wire \output_c[4][19] ;
 wire \output_c[4][1] ;
 wire \output_c[4][20] ;
 wire \output_c[4][21] ;
 wire \output_c[4][22] ;
 wire \output_c[4][23] ;
 wire \output_c[4][24] ;
 wire \output_c[4][25] ;
 wire \output_c[4][26] ;
 wire \output_c[4][27] ;
 wire \output_c[4][28] ;
 wire \output_c[4][29] ;
 wire \output_c[4][2] ;
 wire \output_c[4][30] ;
 wire \output_c[4][31] ;
 wire \output_c[4][3] ;
 wire \output_c[4][4] ;
 wire \output_c[4][5] ;
 wire \output_c[4][6] ;
 wire \output_c[4][7] ;
 wire \output_c[4][8] ;
 wire \output_c[4][9] ;
 wire \output_c[5][0] ;
 wire \output_c[5][10] ;
 wire \output_c[5][11] ;
 wire \output_c[5][12] ;
 wire \output_c[5][13] ;
 wire \output_c[5][14] ;
 wire \output_c[5][15] ;
 wire \output_c[5][16] ;
 wire \output_c[5][17] ;
 wire \output_c[5][18] ;
 wire \output_c[5][19] ;
 wire \output_c[5][1] ;
 wire \output_c[5][20] ;
 wire \output_c[5][21] ;
 wire \output_c[5][22] ;
 wire \output_c[5][23] ;
 wire \output_c[5][24] ;
 wire \output_c[5][25] ;
 wire \output_c[5][26] ;
 wire \output_c[5][27] ;
 wire \output_c[5][28] ;
 wire \output_c[5][29] ;
 wire \output_c[5][2] ;
 wire \output_c[5][30] ;
 wire \output_c[5][31] ;
 wire \output_c[5][3] ;
 wire \output_c[5][4] ;
 wire \output_c[5][5] ;
 wire \output_c[5][6] ;
 wire \output_c[5][7] ;
 wire \output_c[5][8] ;
 wire \output_c[5][9] ;
 wire \output_c[6][0] ;
 wire \output_c[6][10] ;
 wire \output_c[6][11] ;
 wire \output_c[6][12] ;
 wire \output_c[6][13] ;
 wire \output_c[6][14] ;
 wire \output_c[6][15] ;
 wire \output_c[6][16] ;
 wire \output_c[6][17] ;
 wire \output_c[6][18] ;
 wire \output_c[6][19] ;
 wire \output_c[6][1] ;
 wire \output_c[6][20] ;
 wire \output_c[6][21] ;
 wire \output_c[6][22] ;
 wire \output_c[6][23] ;
 wire \output_c[6][24] ;
 wire \output_c[6][25] ;
 wire \output_c[6][26] ;
 wire \output_c[6][27] ;
 wire \output_c[6][28] ;
 wire \output_c[6][29] ;
 wire \output_c[6][2] ;
 wire \output_c[6][30] ;
 wire \output_c[6][31] ;
 wire \output_c[6][3] ;
 wire \output_c[6][4] ;
 wire \output_c[6][5] ;
 wire \output_c[6][6] ;
 wire \output_c[6][7] ;
 wire \output_c[6][8] ;
 wire \output_c[6][9] ;
 wire \output_c[7][0] ;
 wire \output_c[7][10] ;
 wire \output_c[7][11] ;
 wire \output_c[7][12] ;
 wire \output_c[7][13] ;
 wire \output_c[7][14] ;
 wire \output_c[7][15] ;
 wire \output_c[7][16] ;
 wire \output_c[7][17] ;
 wire \output_c[7][18] ;
 wire \output_c[7][19] ;
 wire \output_c[7][1] ;
 wire \output_c[7][20] ;
 wire \output_c[7][21] ;
 wire \output_c[7][22] ;
 wire \output_c[7][23] ;
 wire \output_c[7][24] ;
 wire \output_c[7][25] ;
 wire \output_c[7][26] ;
 wire \output_c[7][27] ;
 wire \output_c[7][28] ;
 wire \output_c[7][29] ;
 wire \output_c[7][2] ;
 wire \output_c[7][30] ;
 wire \output_c[7][31] ;
 wire \output_c[7][3] ;
 wire \output_c[7][4] ;
 wire \output_c[7][5] ;
 wire \output_c[7][6] ;
 wire \output_c[7][7] ;
 wire \output_c[7][8] ;
 wire \output_c[7][9] ;
 wire \output_c[8][0] ;
 wire \output_c[8][10] ;
 wire \output_c[8][11] ;
 wire \output_c[8][12] ;
 wire \output_c[8][13] ;
 wire \output_c[8][14] ;
 wire \output_c[8][15] ;
 wire \output_c[8][16] ;
 wire \output_c[8][17] ;
 wire \output_c[8][18] ;
 wire \output_c[8][19] ;
 wire \output_c[8][1] ;
 wire \output_c[8][20] ;
 wire \output_c[8][21] ;
 wire \output_c[8][22] ;
 wire \output_c[8][23] ;
 wire \output_c[8][24] ;
 wire \output_c[8][25] ;
 wire \output_c[8][26] ;
 wire \output_c[8][27] ;
 wire \output_c[8][28] ;
 wire \output_c[8][29] ;
 wire \output_c[8][2] ;
 wire \output_c[8][30] ;
 wire \output_c[8][31] ;
 wire \output_c[8][3] ;
 wire \output_c[8][4] ;
 wire \output_c[8][5] ;
 wire \output_c[8][6] ;
 wire \output_c[8][7] ;
 wire \output_c[8][8] ;
 wire \output_c[8][9] ;
 wire \output_c[9][0] ;
 wire \output_c[9][10] ;
 wire \output_c[9][11] ;
 wire \output_c[9][12] ;
 wire \output_c[9][13] ;
 wire \output_c[9][14] ;
 wire \output_c[9][15] ;
 wire \output_c[9][16] ;
 wire \output_c[9][17] ;
 wire \output_c[9][18] ;
 wire \output_c[9][19] ;
 wire \output_c[9][1] ;
 wire \output_c[9][20] ;
 wire \output_c[9][21] ;
 wire \output_c[9][22] ;
 wire \output_c[9][23] ;
 wire \output_c[9][24] ;
 wire \output_c[9][25] ;
 wire \output_c[9][26] ;
 wire \output_c[9][27] ;
 wire \output_c[9][28] ;
 wire \output_c[9][29] ;
 wire \output_c[9][2] ;
 wire \output_c[9][30] ;
 wire \output_c[9][31] ;
 wire \output_c[9][3] ;
 wire \output_c[9][4] ;
 wire \output_c[9][5] ;
 wire \output_c[9][6] ;
 wire \output_c[9][7] ;
 wire \output_c[9][8] ;
 wire \output_c[9][9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;

 sky130_fd_sc_hd__and2_1 _2368_ (.A(\output_c[14][27] ),
    .B(\output_c[14][26] ),
    .X(_1066_));
 sky130_fd_sc_hd__and4_1 _2369_ (.A(\output_c[14][15] ),
    .B(\output_c[14][14] ),
    .C(\output_c[14][13] ),
    .D(\output_c[14][12] ),
    .X(_1067_));
 sky130_fd_sc_hd__and4_1 _2370_ (.A(\output_c[14][11] ),
    .B(\output_c[14][10] ),
    .C(\output_c[14][9] ),
    .D(\output_c[14][8] ),
    .X(_1068_));
 sky130_fd_sc_hd__and2_1 _2371_ (.A(_1067_),
    .B(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_2 _2372_ (.A(\input_b[15][0] ),
    .X(_1070_));
 sky130_fd_sc_hd__buf_1 _2373_ (.A(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__and3_1 _2374_ (.A(\output_c[14][0] ),
    .B(_1071_),
    .C(\input_a[14][0] ),
    .X(_1072_));
 sky130_fd_sc_hd__and4_1 _2375_ (.A(\output_c[14][19] ),
    .B(\output_c[14][18] ),
    .C(\output_c[14][17] ),
    .D(\output_c[14][16] ),
    .X(_1073_));
 sky130_fd_sc_hd__and4_1 _2376_ (.A(\output_c[14][7] ),
    .B(\output_c[14][6] ),
    .C(\output_c[14][5] ),
    .D(\output_c[14][4] ),
    .X(_1074_));
 sky130_fd_sc_hd__and3_1 _2377_ (.A(_1072_),
    .B(_1073_),
    .C(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__buf_1 _2378_ (.A(\output_c[14][2] ),
    .X(_1076_));
 sky130_fd_sc_hd__and4_1 _2379_ (.A(\state[1] ),
    .B(\state[0] ),
    .C(\state[2] ),
    .D(\state[3] ),
    .X(_1077_));
 sky130_fd_sc_hd__buf_1 _2380_ (.A(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_2 _2381_ (.A(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__buf_1 _2382_ (.A(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__and4_1 _2383_ (.A(\output_c[14][23] ),
    .B(\output_c[14][22] ),
    .C(\output_c[14][21] ),
    .D(\output_c[14][20] ),
    .X(_1081_));
 sky130_fd_sc_hd__and2_1 _2384_ (.A(\output_c[14][3] ),
    .B(\output_c[14][1] ),
    .X(_1082_));
 sky130_fd_sc_hd__and4_1 _2385_ (.A(_1076_),
    .B(_1080_),
    .C(_1081_),
    .D(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__and4_1 _2386_ (.A(\output_c[14][24] ),
    .B(_1069_),
    .C(_1075_),
    .D(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__and4_1 _2387_ (.A(\output_c[14][28] ),
    .B(\output_c[14][25] ),
    .C(_1066_),
    .D(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__and3_1 _2388_ (.A(\output_c[14][30] ),
    .B(\output_c[14][29] ),
    .C(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__xor2_1 _2389_ (.A(net58),
    .B(_1086_),
    .X(_1065_));
 sky130_fd_sc_hd__a21oi_1 _2390_ (.A1(\output_c[14][29] ),
    .A2(_1085_),
    .B1(net192),
    .Y(_1087_));
 sky130_fd_sc_hd__nor2_1 _2391_ (.A(_1086_),
    .B(net193),
    .Y(_1064_));
 sky130_fd_sc_hd__xor2_1 _2392_ (.A(net267),
    .B(_1085_),
    .X(_1063_));
 sky130_fd_sc_hd__buf_1 _2393_ (.A(_1084_),
    .X(_1088_));
 sky130_fd_sc_hd__a31o_1 _2394_ (.A1(\output_c[14][25] ),
    .A2(_1066_),
    .A3(_1088_),
    .B1(\output_c[14][28] ),
    .X(_1089_));
 sky130_fd_sc_hd__and2b_1 _2395_ (.A_N(_1085_),
    .B(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_1 _2396_ (.A(_1090_),
    .X(_1062_));
 sky130_fd_sc_hd__buf_1 _2397_ (.A(\output_c[14][25] ),
    .X(_1091_));
 sky130_fd_sc_hd__and3_1 _2398_ (.A(\output_c[14][26] ),
    .B(_1091_),
    .C(_1088_),
    .X(_1092_));
 sky130_fd_sc_hd__xor2_1 _2399_ (.A(net104),
    .B(_1092_),
    .X(_1061_));
 sky130_fd_sc_hd__a21oi_1 _2400_ (.A1(_1091_),
    .A2(_1088_),
    .B1(net478),
    .Y(_1093_));
 sky130_fd_sc_hd__nor2_1 _2401_ (.A(_1092_),
    .B(_1093_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand2_1 _2402_ (.A(_1091_),
    .B(_1088_),
    .Y(_1094_));
 sky130_fd_sc_hd__or2_1 _2403_ (.A(\output_c[14][25] ),
    .B(_1084_),
    .X(_1095_));
 sky130_fd_sc_hd__and2_1 _2404_ (.A(_1094_),
    .B(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2405_ (.A(_1096_),
    .X(_1059_));
 sky130_fd_sc_hd__buf_1 _2406_ (.A(_1069_),
    .X(_1097_));
 sky130_fd_sc_hd__and3_1 _2407_ (.A(_1097_),
    .B(_1075_),
    .C(_1083_),
    .X(_1098_));
 sky130_fd_sc_hd__xor2_1 _2408_ (.A(net88),
    .B(_1098_),
    .X(_1058_));
 sky130_fd_sc_hd__buf_1 _2409_ (.A(\output_c[14][21] ),
    .X(_1099_));
 sky130_fd_sc_hd__buf_1 _2410_ (.A(\output_c[14][20] ),
    .X(_1100_));
 sky130_fd_sc_hd__clkbuf_2 _2411_ (.A(_1078_),
    .X(_1101_));
 sky130_fd_sc_hd__and4_1 _2412_ (.A(\output_c[14][1] ),
    .B(\output_c[14][0] ),
    .C(_1071_),
    .D(\input_a[14][0] ),
    .X(_1102_));
 sky130_fd_sc_hd__and4_1 _2413_ (.A(\output_c[14][3] ),
    .B(\output_c[14][2] ),
    .C(_1101_),
    .D(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__and4_1 _2414_ (.A(_1097_),
    .B(_1073_),
    .C(_1074_),
    .D(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__and2_1 _2415_ (.A(_1100_),
    .B(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__and3_1 _2416_ (.A(\output_c[14][22] ),
    .B(_1099_),
    .C(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__xor2_1 _2417_ (.A(net93),
    .B(_1106_),
    .X(_1057_));
 sky130_fd_sc_hd__and3_1 _2418_ (.A(_1099_),
    .B(_1100_),
    .C(_1104_),
    .X(_1107_));
 sky130_fd_sc_hd__xor2_1 _2419_ (.A(net304),
    .B(_1107_),
    .X(_1056_));
 sky130_fd_sc_hd__nor2_1 _2420_ (.A(_1099_),
    .B(_1105_),
    .Y(_1108_));
 sky130_fd_sc_hd__nor2_1 _2421_ (.A(_1107_),
    .B(_1108_),
    .Y(_1055_));
 sky130_fd_sc_hd__nor2_1 _2422_ (.A(_1100_),
    .B(_1104_),
    .Y(_1109_));
 sky130_fd_sc_hd__nor2_1 _2423_ (.A(_1105_),
    .B(_1109_),
    .Y(_1054_));
 sky130_fd_sc_hd__and2_1 _2424_ (.A(_1074_),
    .B(_1103_),
    .X(_1110_));
 sky130_fd_sc_hd__and3_1 _2425_ (.A(\output_c[14][16] ),
    .B(_1097_),
    .C(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__and3_1 _2426_ (.A(\output_c[14][18] ),
    .B(\output_c[14][17] ),
    .C(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__xor2_1 _2427_ (.A(net129),
    .B(_1112_),
    .X(_1053_));
 sky130_fd_sc_hd__buf_1 _2428_ (.A(\output_c[14][17] ),
    .X(_1113_));
 sky130_fd_sc_hd__buf_1 _2429_ (.A(_1111_),
    .X(_1114_));
 sky130_fd_sc_hd__a21oi_1 _2430_ (.A1(_1113_),
    .A2(_1114_),
    .B1(net477),
    .Y(_1115_));
 sky130_fd_sc_hd__nor2_1 _2431_ (.A(_1112_),
    .B(_1115_),
    .Y(_1052_));
 sky130_fd_sc_hd__and2_1 _2432_ (.A(_1113_),
    .B(_1114_),
    .X(_1116_));
 sky130_fd_sc_hd__nor2_1 _2433_ (.A(_1113_),
    .B(_1114_),
    .Y(_1117_));
 sky130_fd_sc_hd__nor2_1 _2434_ (.A(_1116_),
    .B(_1117_),
    .Y(_1051_));
 sky130_fd_sc_hd__buf_1 _2435_ (.A(_1110_),
    .X(_1118_));
 sky130_fd_sc_hd__a21oi_1 _2436_ (.A1(_1097_),
    .A2(_1118_),
    .B1(net434),
    .Y(_1119_));
 sky130_fd_sc_hd__nor2_1 _2437_ (.A(_1114_),
    .B(_1119_),
    .Y(_1050_));
 sky130_fd_sc_hd__and3_1 _2438_ (.A(\output_c[14][12] ),
    .B(_1068_),
    .C(_1110_),
    .X(_1120_));
 sky130_fd_sc_hd__and3_1 _2439_ (.A(\output_c[14][14] ),
    .B(\output_c[14][13] ),
    .C(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__xor2_1 _2440_ (.A(net153),
    .B(_1121_),
    .X(_1049_));
 sky130_fd_sc_hd__buf_1 _2441_ (.A(\output_c[14][13] ),
    .X(_1122_));
 sky130_fd_sc_hd__buf_1 _2442_ (.A(_1120_),
    .X(_1123_));
 sky130_fd_sc_hd__a21oi_1 _2443_ (.A1(_1122_),
    .A2(_1123_),
    .B1(net454),
    .Y(_1124_));
 sky130_fd_sc_hd__nor2_1 _2444_ (.A(_1121_),
    .B(_1124_),
    .Y(_1048_));
 sky130_fd_sc_hd__and2_1 _2445_ (.A(_1122_),
    .B(_1123_),
    .X(_1125_));
 sky130_fd_sc_hd__nor2_1 _2446_ (.A(_1122_),
    .B(_1123_),
    .Y(_1126_));
 sky130_fd_sc_hd__nor2_1 _2447_ (.A(_1125_),
    .B(_1126_),
    .Y(_1047_));
 sky130_fd_sc_hd__a21oi_1 _2448_ (.A1(_1068_),
    .A2(_1118_),
    .B1(net419),
    .Y(_1127_));
 sky130_fd_sc_hd__nor2_1 _2449_ (.A(_1123_),
    .B(_1127_),
    .Y(_1046_));
 sky130_fd_sc_hd__buf_1 _2450_ (.A(\output_c[14][9] ),
    .X(_1128_));
 sky130_fd_sc_hd__and3_1 _2451_ (.A(\output_c[14][8] ),
    .B(_1074_),
    .C(_1103_),
    .X(_1129_));
 sky130_fd_sc_hd__and3_1 _2452_ (.A(\output_c[14][10] ),
    .B(_1128_),
    .C(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__o2bb2a_1 _2453_ (.A1_N(_1068_),
    .A2_N(_1118_),
    .B1(_1130_),
    .B2(net353),
    .X(_1045_));
 sky130_fd_sc_hd__a21o_1 _2454_ (.A1(_1128_),
    .A2(_1129_),
    .B1(\output_c[14][10] ),
    .X(_1131_));
 sky130_fd_sc_hd__and2b_1 _2455_ (.A_N(_1130_),
    .B(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2456_ (.A(_1132_),
    .X(_1044_));
 sky130_fd_sc_hd__xor2_1 _2457_ (.A(_1128_),
    .B(_1129_),
    .X(_1043_));
 sky130_fd_sc_hd__nor2_1 _2458_ (.A(net465),
    .B(_1118_),
    .Y(_1133_));
 sky130_fd_sc_hd__nor2_1 _2459_ (.A(_1129_),
    .B(_1133_),
    .Y(_1042_));
 sky130_fd_sc_hd__buf_1 _2460_ (.A(\output_c[14][5] ),
    .X(_1134_));
 sky130_fd_sc_hd__buf_1 _2461_ (.A(\output_c[14][4] ),
    .X(_1135_));
 sky130_fd_sc_hd__buf_1 _2462_ (.A(_1103_),
    .X(_1136_));
 sky130_fd_sc_hd__and2_1 _2463_ (.A(_1135_),
    .B(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__and3_1 _2464_ (.A(\output_c[14][6] ),
    .B(_1134_),
    .C(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__xor2_1 _2465_ (.A(net91),
    .B(_1138_),
    .X(_1041_));
 sky130_fd_sc_hd__and3_1 _2466_ (.A(_1134_),
    .B(_1135_),
    .C(_1136_),
    .X(_1139_));
 sky130_fd_sc_hd__nor2_1 _2467_ (.A(net464),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__nor2_1 _2468_ (.A(_1138_),
    .B(_1140_),
    .Y(_1040_));
 sky130_fd_sc_hd__nor2_1 _2469_ (.A(_1134_),
    .B(_1137_),
    .Y(_1141_));
 sky130_fd_sc_hd__nor2_1 _2470_ (.A(_1139_),
    .B(_1141_),
    .Y(_1039_));
 sky130_fd_sc_hd__nor2_1 _2471_ (.A(_1135_),
    .B(_1136_),
    .Y(_1142_));
 sky130_fd_sc_hd__nor2_1 _2472_ (.A(_1137_),
    .B(_1142_),
    .Y(_1038_));
 sky130_fd_sc_hd__buf_1 _2473_ (.A(_1080_),
    .X(_1143_));
 sky130_fd_sc_hd__buf_1 _2474_ (.A(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__and3_1 _2475_ (.A(_1076_),
    .B(_1144_),
    .C(_1102_),
    .X(_1145_));
 sky130_fd_sc_hd__nor2_1 _2476_ (.A(net467),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__nor2_1 _2477_ (.A(_1136_),
    .B(_1146_),
    .Y(_1037_));
 sky130_fd_sc_hd__buf_1 _2478_ (.A(_1143_),
    .X(_1147_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2479_ (.A(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__a21oi_1 _2480_ (.A1(_1148_),
    .A2(_1102_),
    .B1(_1076_),
    .Y(_1149_));
 sky130_fd_sc_hd__nor2_1 _2481_ (.A(_1145_),
    .B(_1149_),
    .Y(_1036_));
 sky130_fd_sc_hd__buf_1 _2482_ (.A(_1144_),
    .X(_1150_));
 sky130_fd_sc_hd__a21oi_1 _2483_ (.A1(_1150_),
    .A2(_1072_),
    .B1(net452),
    .Y(_1151_));
 sky130_fd_sc_hd__a21oi_1 _2484_ (.A1(_1148_),
    .A2(_1102_),
    .B1(_1151_),
    .Y(_1035_));
 sky130_fd_sc_hd__buf_1 _2485_ (.A(_1150_),
    .X(_1152_));
 sky130_fd_sc_hd__buf_1 _2486_ (.A(_1071_),
    .X(_1153_));
 sky130_fd_sc_hd__buf_1 _2487_ (.A(_1080_),
    .X(_1154_));
 sky130_fd_sc_hd__buf_1 _2488_ (.A(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__buf_1 _2489_ (.A(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a31o_1 _2490_ (.A1(_1153_),
    .A2(\input_a[14][0] ),
    .A3(_1156_),
    .B1(\output_c[14][0] ),
    .X(_1157_));
 sky130_fd_sc_hd__a21boi_1 _2491_ (.A1(_1152_),
    .A2(_1072_),
    .B1_N(_1157_),
    .Y(_1034_));
 sky130_fd_sc_hd__and4_1 _2492_ (.A(\output_c[13][27] ),
    .B(\output_c[13][26] ),
    .C(\output_c[13][25] ),
    .D(\output_c[13][24] ),
    .X(_1158_));
 sky130_fd_sc_hd__and4_1 _2493_ (.A(\output_c[13][11] ),
    .B(\output_c[13][10] ),
    .C(\output_c[13][9] ),
    .D(\output_c[13][8] ),
    .X(_1159_));
 sky130_fd_sc_hd__and3_1 _2494_ (.A(\output_c[13][13] ),
    .B(\output_c[13][12] ),
    .C(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__and3_1 _2495_ (.A(\output_c[13][15] ),
    .B(\output_c[13][14] ),
    .C(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__buf_1 _2496_ (.A(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__buf_1 _2497_ (.A(\output_c[13][4] ),
    .X(_1163_));
 sky130_fd_sc_hd__clkbuf_2 _2498_ (.A(_1077_),
    .X(_1164_));
 sky130_fd_sc_hd__and3_1 _2499_ (.A(\output_c[13][0] ),
    .B(_1070_),
    .C(\input_a[13][0] ),
    .X(_1165_));
 sky130_fd_sc_hd__and2_1 _2500_ (.A(\output_c[13][3] ),
    .B(\output_c[13][2] ),
    .X(_1166_));
 sky130_fd_sc_hd__and4_1 _2501_ (.A(\output_c[13][1] ),
    .B(_1164_),
    .C(_1165_),
    .D(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__and2_1 _2502_ (.A(\output_c[13][7] ),
    .B(\output_c[13][6] ),
    .X(_1168_));
 sky130_fd_sc_hd__and4_1 _2503_ (.A(\output_c[13][5] ),
    .B(_1163_),
    .C(_1167_),
    .D(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__and2_1 _2504_ (.A(\output_c[13][21] ),
    .B(\output_c[13][20] ),
    .X(_1170_));
 sky130_fd_sc_hd__and4_1 _2505_ (.A(\output_c[13][19] ),
    .B(\output_c[13][18] ),
    .C(\output_c[13][17] ),
    .D(\output_c[13][16] ),
    .X(_1171_));
 sky130_fd_sc_hd__and4_1 _2506_ (.A(\output_c[13][23] ),
    .B(\output_c[13][22] ),
    .C(_1170_),
    .D(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__and4_1 _2507_ (.A(_1158_),
    .B(_1162_),
    .C(_1169_),
    .D(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__and4_1 _2508_ (.A(\output_c[13][30] ),
    .B(\output_c[13][29] ),
    .C(\output_c[13][28] ),
    .D(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__xor2_1 _2509_ (.A(net44),
    .B(_1174_),
    .X(_1033_));
 sky130_fd_sc_hd__and2_1 _2510_ (.A(\output_c[13][6] ),
    .B(\output_c[13][5] ),
    .X(_1175_));
 sky130_fd_sc_hd__and4_1 _2511_ (.A(\output_c[13][7] ),
    .B(\output_c[13][4] ),
    .C(_1167_),
    .D(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__buf_1 _2512_ (.A(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__and4_1 _2513_ (.A(_1158_),
    .B(_1162_),
    .C(_1172_),
    .D(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__and3_1 _2514_ (.A(\output_c[13][29] ),
    .B(\output_c[13][28] ),
    .C(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__xor2_1 _2515_ (.A(net73),
    .B(_1179_),
    .X(_1032_));
 sky130_fd_sc_hd__a21oi_1 _2516_ (.A1(net275),
    .A2(_1178_),
    .B1(net394),
    .Y(_1180_));
 sky130_fd_sc_hd__nor2_1 _2517_ (.A(_1179_),
    .B(_1180_),
    .Y(_1031_));
 sky130_fd_sc_hd__xor2_1 _2518_ (.A(net275),
    .B(_1178_),
    .X(_1030_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2519_ (.A(\output_c[13][24] ),
    .X(_1181_));
 sky130_fd_sc_hd__and3_1 _2520_ (.A(_1161_),
    .B(_1172_),
    .C(_1176_),
    .X(_1182_));
 sky130_fd_sc_hd__a41o_1 _2521_ (.A1(\output_c[13][26] ),
    .A2(\output_c[13][25] ),
    .A3(_1181_),
    .A4(_1182_),
    .B1(\output_c[13][27] ),
    .X(_1183_));
 sky130_fd_sc_hd__and2b_1 _2522_ (.A_N(_1178_),
    .B(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2523_ (.A(_1184_),
    .X(_1029_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2524_ (.A(_1182_),
    .X(_1185_));
 sky130_fd_sc_hd__nand3_1 _2525_ (.A(\output_c[13][25] ),
    .B(_1181_),
    .C(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__xnor2_1 _2526_ (.A(net166),
    .B(_1186_),
    .Y(_1028_));
 sky130_fd_sc_hd__a21o_1 _2527_ (.A1(_1181_),
    .A2(_1185_),
    .B1(\output_c[13][25] ),
    .X(_1187_));
 sky130_fd_sc_hd__and2_1 _2528_ (.A(_1186_),
    .B(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _2529_ (.A(_1188_),
    .X(_1027_));
 sky130_fd_sc_hd__xor2_1 _2530_ (.A(_1181_),
    .B(_1185_),
    .X(_1026_));
 sky130_fd_sc_hd__and4_1 _2531_ (.A(_1162_),
    .B(_1170_),
    .C(_1171_),
    .D(_1177_),
    .X(_1189_));
 sky130_fd_sc_hd__a21oi_1 _2532_ (.A1(\output_c[13][22] ),
    .A2(_1189_),
    .B1(net163),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _2533_ (.A(_1185_),
    .B(net164),
    .Y(_1025_));
 sky130_fd_sc_hd__xor2_1 _2534_ (.A(net176),
    .B(_1189_),
    .X(_1024_));
 sky130_fd_sc_hd__and2_1 _2535_ (.A(_1161_),
    .B(_1177_),
    .X(_1191_));
 sky130_fd_sc_hd__a31o_1 _2536_ (.A1(\output_c[13][20] ),
    .A2(_1171_),
    .A3(_1191_),
    .B1(\output_c[13][21] ),
    .X(_1192_));
 sky130_fd_sc_hd__and2b_1 _2537_ (.A_N(_1189_),
    .B(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2538_ (.A(_1193_),
    .X(_1023_));
 sky130_fd_sc_hd__nand2_1 _2539_ (.A(_1171_),
    .B(_1191_),
    .Y(_1194_));
 sky130_fd_sc_hd__xnor2_1 _2540_ (.A(net236),
    .B(_1194_),
    .Y(_1022_));
 sky130_fd_sc_hd__and3_1 _2541_ (.A(\output_c[13][16] ),
    .B(_1162_),
    .C(_1169_),
    .X(_1195_));
 sky130_fd_sc_hd__and3_1 _2542_ (.A(\output_c[13][18] ),
    .B(\output_c[13][17] ),
    .C(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__o21a_1 _2543_ (.A1(net135),
    .A2(_1196_),
    .B1(_1194_),
    .X(_1021_));
 sky130_fd_sc_hd__a21oi_1 _2544_ (.A1(net297),
    .A2(_1195_),
    .B1(net334),
    .Y(_1197_));
 sky130_fd_sc_hd__nor2_1 _2545_ (.A(_1196_),
    .B(_1197_),
    .Y(_1020_));
 sky130_fd_sc_hd__xor2_1 _2546_ (.A(net297),
    .B(_1195_),
    .X(_1019_));
 sky130_fd_sc_hd__nor2_1 _2547_ (.A(net448),
    .B(_1191_),
    .Y(_1198_));
 sky130_fd_sc_hd__nor2_1 _2548_ (.A(_1195_),
    .B(_1198_),
    .Y(_1018_));
 sky130_fd_sc_hd__and3_1 _2549_ (.A(\output_c[13][12] ),
    .B(_1159_),
    .C(_1169_),
    .X(_1199_));
 sky130_fd_sc_hd__and3_1 _2550_ (.A(\output_c[13][14] ),
    .B(\output_c[13][13] ),
    .C(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__xor2_1 _2551_ (.A(net63),
    .B(_1200_),
    .X(_1017_));
 sky130_fd_sc_hd__buf_1 _2552_ (.A(_1177_),
    .X(_1201_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2553_ (.A(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__a21oi_1 _2554_ (.A1(_1160_),
    .A2(_1202_),
    .B1(net294),
    .Y(_1203_));
 sky130_fd_sc_hd__nor2_1 _2555_ (.A(_1200_),
    .B(_1203_),
    .Y(_1016_));
 sky130_fd_sc_hd__nor2_1 _2556_ (.A(net279),
    .B(_1199_),
    .Y(_1204_));
 sky130_fd_sc_hd__a21oi_1 _2557_ (.A1(_1160_),
    .A2(_1202_),
    .B1(_1204_),
    .Y(_1015_));
 sky130_fd_sc_hd__and2_1 _2558_ (.A(_1159_),
    .B(_1201_),
    .X(_1205_));
 sky130_fd_sc_hd__nor2_1 _2559_ (.A(net391),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__nor2_1 _2560_ (.A(_1199_),
    .B(_1206_),
    .Y(_1014_));
 sky130_fd_sc_hd__and3_1 _2561_ (.A(\output_c[13][9] ),
    .B(\output_c[13][8] ),
    .C(_1201_),
    .X(_1207_));
 sky130_fd_sc_hd__a21oi_1 _2562_ (.A1(\output_c[13][10] ),
    .A2(_1207_),
    .B1(net98),
    .Y(_1208_));
 sky130_fd_sc_hd__nor2_1 _2563_ (.A(_1205_),
    .B(net99),
    .Y(_1013_));
 sky130_fd_sc_hd__xor2_1 _2564_ (.A(net178),
    .B(_1207_),
    .X(_1012_));
 sky130_fd_sc_hd__a21oi_1 _2565_ (.A1(net339),
    .A2(_1202_),
    .B1(net383),
    .Y(_1209_));
 sky130_fd_sc_hd__nor2_1 _2566_ (.A(_1207_),
    .B(_1209_),
    .Y(_1011_));
 sky130_fd_sc_hd__xor2_1 _2567_ (.A(net339),
    .B(_1202_),
    .X(_1010_));
 sky130_fd_sc_hd__buf_1 _2568_ (.A(_1167_),
    .X(_1210_));
 sky130_fd_sc_hd__and3_1 _2569_ (.A(\output_c[13][5] ),
    .B(_1163_),
    .C(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__a21o_1 _2570_ (.A1(\output_c[13][6] ),
    .A2(_1211_),
    .B1(\output_c[13][7] ),
    .X(_1212_));
 sky130_fd_sc_hd__and2b_1 _2571_ (.A_N(_1201_),
    .B(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_1 _2572_ (.A(_1213_),
    .X(_1009_));
 sky130_fd_sc_hd__xor2_1 _2573_ (.A(net268),
    .B(_1211_),
    .X(_1008_));
 sky130_fd_sc_hd__a21oi_1 _2574_ (.A1(_1163_),
    .A2(_1210_),
    .B1(net461),
    .Y(_1214_));
 sky130_fd_sc_hd__nor2_1 _2575_ (.A(_1211_),
    .B(_1214_),
    .Y(_1007_));
 sky130_fd_sc_hd__xor2_1 _2576_ (.A(_1163_),
    .B(_1210_),
    .X(_1006_));
 sky130_fd_sc_hd__buf_1 _2577_ (.A(_1080_),
    .X(_1215_));
 sky130_fd_sc_hd__and3_1 _2578_ (.A(\output_c[13][1] ),
    .B(_1215_),
    .C(_1165_),
    .X(_1216_));
 sky130_fd_sc_hd__and2_1 _2579_ (.A(\output_c[13][2] ),
    .B(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__o21ba_1 _2580_ (.A1(net395),
    .A2(_1217_),
    .B1_N(_1210_),
    .X(_1005_));
 sky130_fd_sc_hd__nor2_1 _2581_ (.A(net418),
    .B(_1216_),
    .Y(_1218_));
 sky130_fd_sc_hd__nor2_1 _2582_ (.A(_1217_),
    .B(_1218_),
    .Y(_1004_));
 sky130_fd_sc_hd__a21oi_1 _2583_ (.A1(_1148_),
    .A2(_1165_),
    .B1(net396),
    .Y(_1219_));
 sky130_fd_sc_hd__nor2_1 _2584_ (.A(_1216_),
    .B(_1219_),
    .Y(_1003_));
 sky130_fd_sc_hd__buf_1 _2585_ (.A(_1215_),
    .X(_1220_));
 sky130_fd_sc_hd__and3_1 _2586_ (.A(_1153_),
    .B(\input_a[13][0] ),
    .C(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__o2bb2a_1 _2587_ (.A1_N(_1152_),
    .A2_N(_1165_),
    .B1(_1221_),
    .B2(net194),
    .X(_1002_));
 sky130_fd_sc_hd__and4_1 _2588_ (.A(\output_c[12][27] ),
    .B(\output_c[12][26] ),
    .C(\output_c[12][25] ),
    .D(\output_c[12][24] ),
    .X(_1222_));
 sky130_fd_sc_hd__and4_1 _2589_ (.A(\output_c[12][11] ),
    .B(\output_c[12][10] ),
    .C(\output_c[12][9] ),
    .D(\output_c[12][8] ),
    .X(_1223_));
 sky130_fd_sc_hd__and3_1 _2590_ (.A(\output_c[12][13] ),
    .B(\output_c[12][12] ),
    .C(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__and3_1 _2591_ (.A(\output_c[12][15] ),
    .B(\output_c[12][14] ),
    .C(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__buf_1 _2592_ (.A(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__buf_1 _2593_ (.A(\output_c[12][4] ),
    .X(_1227_));
 sky130_fd_sc_hd__and3_1 _2594_ (.A(\output_c[12][0] ),
    .B(_1070_),
    .C(\input_a[12][0] ),
    .X(_1228_));
 sky130_fd_sc_hd__and2_1 _2595_ (.A(\output_c[12][3] ),
    .B(\output_c[12][2] ),
    .X(_1229_));
 sky130_fd_sc_hd__and4_1 _2596_ (.A(\output_c[12][1] ),
    .B(_1078_),
    .C(_1228_),
    .D(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__and2_1 _2597_ (.A(\output_c[12][7] ),
    .B(\output_c[12][6] ),
    .X(_1231_));
 sky130_fd_sc_hd__and4_1 _2598_ (.A(\output_c[12][5] ),
    .B(_1227_),
    .C(_1230_),
    .D(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__and2_1 _2599_ (.A(\output_c[12][21] ),
    .B(\output_c[12][20] ),
    .X(_1233_));
 sky130_fd_sc_hd__and4_1 _2600_ (.A(\output_c[12][19] ),
    .B(\output_c[12][18] ),
    .C(\output_c[12][17] ),
    .D(\output_c[12][16] ),
    .X(_1234_));
 sky130_fd_sc_hd__and4_1 _2601_ (.A(\output_c[12][23] ),
    .B(\output_c[12][22] ),
    .C(_1233_),
    .D(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__and4_1 _2602_ (.A(_1222_),
    .B(_1226_),
    .C(_1232_),
    .D(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__and4_1 _2603_ (.A(net495),
    .B(\output_c[12][29] ),
    .C(\output_c[12][28] ),
    .D(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__xor2_1 _2604_ (.A(net41),
    .B(_1237_),
    .X(_1001_));
 sky130_fd_sc_hd__and2_1 _2605_ (.A(\output_c[12][6] ),
    .B(\output_c[12][5] ),
    .X(_1238_));
 sky130_fd_sc_hd__and4_1 _2606_ (.A(\output_c[12][7] ),
    .B(\output_c[12][4] ),
    .C(_1230_),
    .D(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__buf_1 _2607_ (.A(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__and4_1 _2608_ (.A(_1222_),
    .B(_1226_),
    .C(_1235_),
    .D(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__and3_1 _2609_ (.A(\output_c[12][29] ),
    .B(\output_c[12][28] ),
    .C(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__xor2_1 _2610_ (.A(net62),
    .B(_1242_),
    .X(_1000_));
 sky130_fd_sc_hd__a21oi_1 _2611_ (.A1(net296),
    .A2(_1241_),
    .B1(net380),
    .Y(_1243_));
 sky130_fd_sc_hd__nor2_1 _2612_ (.A(_1242_),
    .B(_1243_),
    .Y(_0999_));
 sky130_fd_sc_hd__xor2_1 _2613_ (.A(net296),
    .B(_1241_),
    .X(_0998_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2614_ (.A(\output_c[12][24] ),
    .X(_1244_));
 sky130_fd_sc_hd__and3_1 _2615_ (.A(_1225_),
    .B(_1235_),
    .C(_1239_),
    .X(_1245_));
 sky130_fd_sc_hd__a41o_1 _2616_ (.A1(\output_c[12][26] ),
    .A2(\output_c[12][25] ),
    .A3(_1244_),
    .A4(_1245_),
    .B1(\output_c[12][27] ),
    .X(_1246_));
 sky130_fd_sc_hd__and2b_1 _2617_ (.A_N(_1241_),
    .B(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _2618_ (.A(_1247_),
    .X(_0997_));
 sky130_fd_sc_hd__buf_1 _2619_ (.A(_1245_),
    .X(_1248_));
 sky130_fd_sc_hd__nand3_1 _2620_ (.A(\output_c[12][25] ),
    .B(_1244_),
    .C(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__xnor2_1 _2621_ (.A(net186),
    .B(_1249_),
    .Y(_0996_));
 sky130_fd_sc_hd__a21o_1 _2622_ (.A1(_1244_),
    .A2(_1248_),
    .B1(\output_c[12][25] ),
    .X(_1250_));
 sky130_fd_sc_hd__and2_1 _2623_ (.A(_1249_),
    .B(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _2624_ (.A(_1251_),
    .X(_0995_));
 sky130_fd_sc_hd__xor2_1 _2625_ (.A(_1244_),
    .B(_1248_),
    .X(_0994_));
 sky130_fd_sc_hd__and4_1 _2626_ (.A(_1226_),
    .B(_1233_),
    .C(_1234_),
    .D(_1240_),
    .X(_1252_));
 sky130_fd_sc_hd__a21oi_1 _2627_ (.A1(\output_c[12][22] ),
    .A2(_1252_),
    .B1(net149),
    .Y(_1253_));
 sky130_fd_sc_hd__nor2_1 _2628_ (.A(_1248_),
    .B(net150),
    .Y(_0993_));
 sky130_fd_sc_hd__xor2_1 _2629_ (.A(net172),
    .B(_1252_),
    .X(_0992_));
 sky130_fd_sc_hd__and2_1 _2630_ (.A(_1225_),
    .B(_1240_),
    .X(_1254_));
 sky130_fd_sc_hd__a31o_1 _2631_ (.A1(\output_c[12][20] ),
    .A2(_1234_),
    .A3(_1254_),
    .B1(\output_c[12][21] ),
    .X(_1255_));
 sky130_fd_sc_hd__and2b_1 _2632_ (.A_N(_1252_),
    .B(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_1256_),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_1 _2634_ (.A(_1234_),
    .B(_1254_),
    .Y(_1257_));
 sky130_fd_sc_hd__xnor2_1 _2635_ (.A(net130),
    .B(_1257_),
    .Y(_0990_));
 sky130_fd_sc_hd__and3_1 _2636_ (.A(\output_c[12][16] ),
    .B(_1226_),
    .C(_1232_),
    .X(_1258_));
 sky130_fd_sc_hd__and3_1 _2637_ (.A(\output_c[12][18] ),
    .B(\output_c[12][17] ),
    .C(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__o21a_1 _2638_ (.A1(net87),
    .A2(_1259_),
    .B1(_1257_),
    .X(_0989_));
 sky130_fd_sc_hd__a21oi_1 _2639_ (.A1(\output_c[12][17] ),
    .A2(_1258_),
    .B1(net214),
    .Y(_1260_));
 sky130_fd_sc_hd__nor2_1 _2640_ (.A(_1259_),
    .B(net215),
    .Y(_0988_));
 sky130_fd_sc_hd__xor2_1 _2641_ (.A(net269),
    .B(_1258_),
    .X(_0987_));
 sky130_fd_sc_hd__nor2_1 _2642_ (.A(net326),
    .B(_1254_),
    .Y(_1261_));
 sky130_fd_sc_hd__nor2_1 _2643_ (.A(_1258_),
    .B(_1261_),
    .Y(_0986_));
 sky130_fd_sc_hd__and3_1 _2644_ (.A(\output_c[12][12] ),
    .B(_1223_),
    .C(_1232_),
    .X(_1262_));
 sky130_fd_sc_hd__and3_1 _2645_ (.A(\output_c[12][14] ),
    .B(net201),
    .C(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__xor2_1 _2646_ (.A(net53),
    .B(_1263_),
    .X(_0985_));
 sky130_fd_sc_hd__buf_1 _2647_ (.A(_1240_),
    .X(_1264_));
 sky130_fd_sc_hd__buf_1 _2648_ (.A(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__a21oi_1 _2649_ (.A1(_1224_),
    .A2(_1265_),
    .B1(net458),
    .Y(_1266_));
 sky130_fd_sc_hd__nor2_1 _2650_ (.A(_1263_),
    .B(_1266_),
    .Y(_0984_));
 sky130_fd_sc_hd__nor2_1 _2651_ (.A(net201),
    .B(_1262_),
    .Y(_1267_));
 sky130_fd_sc_hd__a21oi_1 _2652_ (.A1(_1224_),
    .A2(_1265_),
    .B1(_1267_),
    .Y(_0983_));
 sky130_fd_sc_hd__and2_1 _2653_ (.A(_1223_),
    .B(_1264_),
    .X(_1268_));
 sky130_fd_sc_hd__nor2_1 _2654_ (.A(net369),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__nor2_1 _2655_ (.A(_1262_),
    .B(_1269_),
    .Y(_0982_));
 sky130_fd_sc_hd__and3_1 _2656_ (.A(\output_c[12][9] ),
    .B(\output_c[12][8] ),
    .C(_1264_),
    .X(_1270_));
 sky130_fd_sc_hd__a21oi_1 _2657_ (.A1(net138),
    .A2(_1270_),
    .B1(net143),
    .Y(_1271_));
 sky130_fd_sc_hd__nor2_1 _2658_ (.A(_1268_),
    .B(_1271_),
    .Y(_0981_));
 sky130_fd_sc_hd__xor2_1 _2659_ (.A(net138),
    .B(_1270_),
    .X(_0980_));
 sky130_fd_sc_hd__a21oi_1 _2660_ (.A1(net308),
    .A2(_1265_),
    .B1(net313),
    .Y(_1272_));
 sky130_fd_sc_hd__nor2_1 _2661_ (.A(_1270_),
    .B(_1272_),
    .Y(_0979_));
 sky130_fd_sc_hd__xor2_1 _2662_ (.A(net308),
    .B(_1265_),
    .X(_0978_));
 sky130_fd_sc_hd__buf_1 _2663_ (.A(_1230_),
    .X(_1273_));
 sky130_fd_sc_hd__and3_1 _2664_ (.A(\output_c[12][5] ),
    .B(_1227_),
    .C(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a21o_1 _2665_ (.A1(\output_c[12][6] ),
    .A2(_1274_),
    .B1(\output_c[12][7] ),
    .X(_1275_));
 sky130_fd_sc_hd__and2b_1 _2666_ (.A_N(_1264_),
    .B(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _2667_ (.A(_1276_),
    .X(_0977_));
 sky130_fd_sc_hd__xor2_1 _2668_ (.A(net309),
    .B(_1274_),
    .X(_0976_));
 sky130_fd_sc_hd__a21oi_1 _2669_ (.A1(_1227_),
    .A2(_1273_),
    .B1(net449),
    .Y(_1277_));
 sky130_fd_sc_hd__nor2_1 _2670_ (.A(_1274_),
    .B(_1277_),
    .Y(_0975_));
 sky130_fd_sc_hd__xor2_1 _2671_ (.A(_1227_),
    .B(_1273_),
    .X(_0974_));
 sky130_fd_sc_hd__and3_1 _2672_ (.A(\output_c[12][1] ),
    .B(_1215_),
    .C(_1228_),
    .X(_1278_));
 sky130_fd_sc_hd__and2_1 _2673_ (.A(net408),
    .B(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__o21ba_1 _2674_ (.A1(net264),
    .A2(_1279_),
    .B1_N(_1273_),
    .X(_0973_));
 sky130_fd_sc_hd__nor2_1 _2675_ (.A(net408),
    .B(_1278_),
    .Y(_1280_));
 sky130_fd_sc_hd__nor2_1 _2676_ (.A(_1279_),
    .B(_1280_),
    .Y(_0972_));
 sky130_fd_sc_hd__a21oi_1 _2677_ (.A1(_1148_),
    .A2(_1228_),
    .B1(net283),
    .Y(_1281_));
 sky130_fd_sc_hd__nor2_1 _2678_ (.A(_1278_),
    .B(_1281_),
    .Y(_0971_));
 sky130_fd_sc_hd__and3_1 _2679_ (.A(_1153_),
    .B(\input_a[12][0] ),
    .C(_1220_),
    .X(_1282_));
 sky130_fd_sc_hd__o2bb2a_1 _2680_ (.A1_N(_1152_),
    .A2_N(_1228_),
    .B1(_1282_),
    .B2(net173),
    .X(_0970_));
 sky130_fd_sc_hd__and4_1 _2681_ (.A(\output_c[11][27] ),
    .B(\output_c[11][26] ),
    .C(\output_c[11][25] ),
    .D(\output_c[11][24] ),
    .X(_1283_));
 sky130_fd_sc_hd__and4_1 _2682_ (.A(\output_c[11][11] ),
    .B(\output_c[11][10] ),
    .C(\output_c[11][9] ),
    .D(\output_c[11][8] ),
    .X(_1284_));
 sky130_fd_sc_hd__and3_1 _2683_ (.A(\output_c[11][13] ),
    .B(\output_c[11][12] ),
    .C(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__and3_1 _2684_ (.A(\output_c[11][15] ),
    .B(\output_c[11][14] ),
    .C(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__buf_1 _2685_ (.A(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_2 _2686_ (.A(_1078_),
    .X(_1288_));
 sky130_fd_sc_hd__buf_1 _2687_ (.A(\input_b[15][0] ),
    .X(_1289_));
 sky130_fd_sc_hd__and3_1 _2688_ (.A(\output_c[11][0] ),
    .B(_1289_),
    .C(\input_a[11][0] ),
    .X(_1290_));
 sky130_fd_sc_hd__and2_1 _2689_ (.A(\output_c[11][3] ),
    .B(\output_c[11][2] ),
    .X(_1291_));
 sky130_fd_sc_hd__and4_1 _2690_ (.A(\output_c[11][1] ),
    .B(_1288_),
    .C(_1290_),
    .D(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__and2_1 _2691_ (.A(\output_c[11][7] ),
    .B(\output_c[11][6] ),
    .X(_1293_));
 sky130_fd_sc_hd__and4_1 _2692_ (.A(\output_c[11][5] ),
    .B(\output_c[11][4] ),
    .C(_1292_),
    .D(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__buf_1 _2693_ (.A(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__and2_1 _2694_ (.A(\output_c[11][21] ),
    .B(\output_c[11][20] ),
    .X(_1296_));
 sky130_fd_sc_hd__and4_1 _2695_ (.A(\output_c[11][19] ),
    .B(\output_c[11][18] ),
    .C(\output_c[11][17] ),
    .D(\output_c[11][16] ),
    .X(_1297_));
 sky130_fd_sc_hd__and2_1 _2696_ (.A(_1296_),
    .B(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__and3_1 _2697_ (.A(\output_c[11][23] ),
    .B(\output_c[11][22] ),
    .C(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__and4_1 _2698_ (.A(_1283_),
    .B(_1287_),
    .C(_1295_),
    .D(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__and4_1 _2699_ (.A(\output_c[11][30] ),
    .B(\output_c[11][29] ),
    .C(\output_c[11][28] ),
    .D(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__xor2_1 _2700_ (.A(net39),
    .B(_1301_),
    .X(_0969_));
 sky130_fd_sc_hd__buf_1 _2701_ (.A(\output_c[11][4] ),
    .X(_1302_));
 sky130_fd_sc_hd__and2_1 _2702_ (.A(\output_c[11][6] ),
    .B(\output_c[11][5] ),
    .X(_1303_));
 sky130_fd_sc_hd__and4_1 _2703_ (.A(\output_c[11][7] ),
    .B(_1302_),
    .C(_1292_),
    .D(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__buf_1 _2704_ (.A(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__and4_1 _2705_ (.A(\output_c[11][23] ),
    .B(\output_c[11][22] ),
    .C(_1296_),
    .D(_1297_),
    .X(_1306_));
 sky130_fd_sc_hd__and3_1 _2706_ (.A(_1287_),
    .B(_1305_),
    .C(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__and4_1 _2707_ (.A(\output_c[11][29] ),
    .B(\output_c[11][28] ),
    .C(_1283_),
    .D(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__xor2_1 _2708_ (.A(net72),
    .B(_1308_),
    .X(_0968_));
 sky130_fd_sc_hd__a21oi_1 _2709_ (.A1(net336),
    .A2(_1300_),
    .B1(net385),
    .Y(_1309_));
 sky130_fd_sc_hd__nor2_1 _2710_ (.A(_1308_),
    .B(_1309_),
    .Y(_0967_));
 sky130_fd_sc_hd__xor2_1 _2711_ (.A(net336),
    .B(_1300_),
    .X(_0966_));
 sky130_fd_sc_hd__buf_1 _2712_ (.A(_1286_),
    .X(_1310_));
 sky130_fd_sc_hd__and4_1 _2713_ (.A(\output_c[11][24] ),
    .B(_1310_),
    .C(_1295_),
    .D(_1299_),
    .X(_1311_));
 sky130_fd_sc_hd__and3_1 _2714_ (.A(\output_c[11][26] ),
    .B(\output_c[11][25] ),
    .C(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__o21ba_1 _2715_ (.A1(net126),
    .A2(_1312_),
    .B1_N(_1300_),
    .X(_0965_));
 sky130_fd_sc_hd__nand2_1 _2716_ (.A(net492),
    .B(_1311_),
    .Y(_1313_));
 sky130_fd_sc_hd__xnor2_1 _2717_ (.A(net97),
    .B(_1313_),
    .Y(_0964_));
 sky130_fd_sc_hd__xor2_1 _2718_ (.A(net370),
    .B(_1311_),
    .X(_0963_));
 sky130_fd_sc_hd__nor2_1 _2719_ (.A(net349),
    .B(_1307_),
    .Y(_1314_));
 sky130_fd_sc_hd__nor2_1 _2720_ (.A(_1311_),
    .B(_1314_),
    .Y(_0962_));
 sky130_fd_sc_hd__and4_1 _2721_ (.A(\output_c[11][22] ),
    .B(_1310_),
    .C(_1295_),
    .D(_1298_),
    .X(_1315_));
 sky130_fd_sc_hd__xor2_1 _2722_ (.A(net89),
    .B(_1315_),
    .X(_0961_));
 sky130_fd_sc_hd__and3_1 _2723_ (.A(_1287_),
    .B(_1297_),
    .C(_1304_),
    .X(_1316_));
 sky130_fd_sc_hd__nand2_1 _2724_ (.A(_1296_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__xnor2_1 _2725_ (.A(net293),
    .B(_1317_),
    .Y(_0960_));
 sky130_fd_sc_hd__a21o_1 _2726_ (.A1(\output_c[11][20] ),
    .A2(_1316_),
    .B1(\output_c[11][21] ),
    .X(_1318_));
 sky130_fd_sc_hd__and2_1 _2727_ (.A(_1317_),
    .B(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _2728_ (.A(_1319_),
    .X(_0959_));
 sky130_fd_sc_hd__xor2_1 _2729_ (.A(net154),
    .B(_1316_),
    .X(_0958_));
 sky130_fd_sc_hd__and4_1 _2730_ (.A(\output_c[11][17] ),
    .B(\output_c[11][16] ),
    .C(_1287_),
    .D(_1294_),
    .X(_1320_));
 sky130_fd_sc_hd__a21o_1 _2731_ (.A1(\output_c[11][18] ),
    .A2(_1320_),
    .B1(\output_c[11][19] ),
    .X(_1321_));
 sky130_fd_sc_hd__and2b_1 _2732_ (.A_N(_1316_),
    .B(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _2733_ (.A(_1322_),
    .X(_0957_));
 sky130_fd_sc_hd__xor2_1 _2734_ (.A(net132),
    .B(_1320_),
    .X(_0956_));
 sky130_fd_sc_hd__and3_1 _2735_ (.A(\output_c[11][16] ),
    .B(_1310_),
    .C(_1305_),
    .X(_1323_));
 sky130_fd_sc_hd__nor2_1 _2736_ (.A(net374),
    .B(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__nor2_1 _2737_ (.A(_1320_),
    .B(_1324_),
    .Y(_0955_));
 sky130_fd_sc_hd__buf_1 _2738_ (.A(_1305_),
    .X(_1325_));
 sky130_fd_sc_hd__buf_1 _2739_ (.A(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__a21oi_1 _2740_ (.A1(_1310_),
    .A2(_1326_),
    .B1(net401),
    .Y(_1327_));
 sky130_fd_sc_hd__nor2_1 _2741_ (.A(_1323_),
    .B(_1327_),
    .Y(_0954_));
 sky130_fd_sc_hd__and3_1 _2742_ (.A(\output_c[11][12] ),
    .B(_1284_),
    .C(_1295_),
    .X(_1328_));
 sky130_fd_sc_hd__and3_1 _2743_ (.A(\output_c[11][14] ),
    .B(\output_c[11][13] ),
    .C(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__xor2_1 _2744_ (.A(net71),
    .B(_1329_),
    .X(_0953_));
 sky130_fd_sc_hd__a21oi_1 _2745_ (.A1(_1285_),
    .A2(_1326_),
    .B1(net288),
    .Y(_1330_));
 sky130_fd_sc_hd__nor2_1 _2746_ (.A(_1329_),
    .B(_1330_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2_1 _2747_ (.A(net232),
    .B(_1328_),
    .Y(_1331_));
 sky130_fd_sc_hd__a21oi_1 _2748_ (.A1(_1285_),
    .A2(_1326_),
    .B1(_1331_),
    .Y(_0951_));
 sky130_fd_sc_hd__and2_1 _2749_ (.A(_1284_),
    .B(_1325_),
    .X(_1332_));
 sky130_fd_sc_hd__nor2_1 _2750_ (.A(net441),
    .B(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__nor2_1 _2751_ (.A(_1328_),
    .B(_1333_),
    .Y(_0950_));
 sky130_fd_sc_hd__and3_1 _2752_ (.A(\output_c[11][9] ),
    .B(\output_c[11][8] ),
    .C(_1305_),
    .X(_1334_));
 sky130_fd_sc_hd__a21oi_1 _2753_ (.A1(\output_c[11][10] ),
    .A2(_1334_),
    .B1(net112),
    .Y(_1335_));
 sky130_fd_sc_hd__nor2_1 _2754_ (.A(_1332_),
    .B(net113),
    .Y(_0949_));
 sky130_fd_sc_hd__xor2_1 _2755_ (.A(net159),
    .B(_1334_),
    .X(_0948_));
 sky130_fd_sc_hd__a21oi_1 _2756_ (.A1(net328),
    .A2(_1325_),
    .B1(net411),
    .Y(_1336_));
 sky130_fd_sc_hd__nor2_1 _2757_ (.A(_1334_),
    .B(_1336_),
    .Y(_0947_));
 sky130_fd_sc_hd__xor2_1 _2758_ (.A(net328),
    .B(_1326_),
    .X(_0946_));
 sky130_fd_sc_hd__buf_1 _2759_ (.A(_1292_),
    .X(_1337_));
 sky130_fd_sc_hd__and3_1 _2760_ (.A(\output_c[11][5] ),
    .B(_1302_),
    .C(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__a21o_1 _2761_ (.A1(\output_c[11][6] ),
    .A2(_1338_),
    .B1(\output_c[11][7] ),
    .X(_1339_));
 sky130_fd_sc_hd__and2b_1 _2762_ (.A_N(_1325_),
    .B(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _2763_ (.A(_1340_),
    .X(_0945_));
 sky130_fd_sc_hd__xor2_1 _2764_ (.A(net335),
    .B(_1338_),
    .X(_0944_));
 sky130_fd_sc_hd__a21oi_1 _2765_ (.A1(_1302_),
    .A2(_1337_),
    .B1(net460),
    .Y(_1341_));
 sky130_fd_sc_hd__nor2_1 _2766_ (.A(_1338_),
    .B(_1341_),
    .Y(_0943_));
 sky130_fd_sc_hd__xor2_1 _2767_ (.A(_1302_),
    .B(_1337_),
    .X(_0942_));
 sky130_fd_sc_hd__and3_1 _2768_ (.A(\output_c[11][1] ),
    .B(_1215_),
    .C(_1290_),
    .X(_1342_));
 sky130_fd_sc_hd__and2_1 _2769_ (.A(\output_c[11][2] ),
    .B(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__o21ba_1 _2770_ (.A1(net227),
    .A2(_1343_),
    .B1_N(_1337_),
    .X(_0941_));
 sky130_fd_sc_hd__nor2_1 _2771_ (.A(net424),
    .B(_1342_),
    .Y(_1344_));
 sky130_fd_sc_hd__nor2_1 _2772_ (.A(_1343_),
    .B(_1344_),
    .Y(_0940_));
 sky130_fd_sc_hd__buf_1 _2773_ (.A(_1143_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_2 _2774_ (.A(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a21oi_1 _2775_ (.A1(_1346_),
    .A2(_1290_),
    .B1(net381),
    .Y(_1347_));
 sky130_fd_sc_hd__nor2_1 _2776_ (.A(_1342_),
    .B(_1347_),
    .Y(_0939_));
 sky130_fd_sc_hd__buf_1 _2777_ (.A(_1071_),
    .X(_1348_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2778_ (.A(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__and3_1 _2779_ (.A(_1349_),
    .B(\input_a[11][0] ),
    .C(_1220_),
    .X(_1350_));
 sky130_fd_sc_hd__o2bb2a_1 _2780_ (.A1_N(_1152_),
    .A2_N(_1290_),
    .B1(_1350_),
    .B2(net142),
    .X(_0938_));
 sky130_fd_sc_hd__and4_1 _2781_ (.A(\output_c[10][27] ),
    .B(\output_c[10][26] ),
    .C(\output_c[10][25] ),
    .D(\output_c[10][24] ),
    .X(_1351_));
 sky130_fd_sc_hd__and4_1 _2782_ (.A(\output_c[10][19] ),
    .B(\output_c[10][18] ),
    .C(\output_c[10][17] ),
    .D(\output_c[10][16] ),
    .X(_1352_));
 sky130_fd_sc_hd__and3_1 _2783_ (.A(\output_c[10][21] ),
    .B(\output_c[10][20] ),
    .C(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__and3_1 _2784_ (.A(\output_c[10][23] ),
    .B(\output_c[10][22] ),
    .C(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__buf_1 _2785_ (.A(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__and4_1 _2786_ (.A(\output_c[10][11] ),
    .B(\output_c[10][10] ),
    .C(\output_c[10][9] ),
    .D(\output_c[10][8] ),
    .X(_1356_));
 sky130_fd_sc_hd__and3_1 _2787_ (.A(\output_c[10][13] ),
    .B(net295),
    .C(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__and3_1 _2788_ (.A(\output_c[10][15] ),
    .B(\output_c[10][14] ),
    .C(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__buf_1 _2789_ (.A(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__buf_1 _2790_ (.A(\output_c[10][4] ),
    .X(_1360_));
 sky130_fd_sc_hd__and3_1 _2791_ (.A(\output_c[10][0] ),
    .B(_1289_),
    .C(\input_a[10][0] ),
    .X(_1361_));
 sky130_fd_sc_hd__and2_1 _2792_ (.A(\output_c[10][3] ),
    .B(\output_c[10][2] ),
    .X(_1362_));
 sky130_fd_sc_hd__and4_1 _2793_ (.A(\output_c[10][1] ),
    .B(_1164_),
    .C(_1361_),
    .D(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__and2_1 _2794_ (.A(\output_c[10][7] ),
    .B(\output_c[10][6] ),
    .X(_1364_));
 sky130_fd_sc_hd__and4_1 _2795_ (.A(\output_c[10][5] ),
    .B(_1360_),
    .C(_1363_),
    .D(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__and4_1 _2796_ (.A(_1351_),
    .B(_1355_),
    .C(_1359_),
    .D(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__and4_1 _2797_ (.A(net493),
    .B(\output_c[10][29] ),
    .C(\output_c[10][28] ),
    .D(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__xor2_1 _2798_ (.A(net37),
    .B(_1367_),
    .X(_0937_));
 sky130_fd_sc_hd__and2_1 _2799_ (.A(\output_c[10][6] ),
    .B(\output_c[10][5] ),
    .X(_1368_));
 sky130_fd_sc_hd__and4_1 _2800_ (.A(\output_c[10][7] ),
    .B(\output_c[10][4] ),
    .C(_1363_),
    .D(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__buf_1 _2801_ (.A(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__and4_1 _2802_ (.A(_1351_),
    .B(_1355_),
    .C(_1359_),
    .D(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__and3_1 _2803_ (.A(\output_c[10][29] ),
    .B(\output_c[10][28] ),
    .C(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__xor2_1 _2804_ (.A(net70),
    .B(_1372_),
    .X(_0936_));
 sky130_fd_sc_hd__a21oi_1 _2805_ (.A1(net260),
    .A2(_1371_),
    .B1(net321),
    .Y(_1373_));
 sky130_fd_sc_hd__nor2_1 _2806_ (.A(_1372_),
    .B(_1373_),
    .Y(_0935_));
 sky130_fd_sc_hd__xor2_1 _2807_ (.A(net260),
    .B(_1371_),
    .X(_0934_));
 sky130_fd_sc_hd__buf_1 _2808_ (.A(\output_c[10][24] ),
    .X(_1374_));
 sky130_fd_sc_hd__and3_1 _2809_ (.A(_1354_),
    .B(_1358_),
    .C(_1369_),
    .X(_1375_));
 sky130_fd_sc_hd__a41o_1 _2810_ (.A1(\output_c[10][26] ),
    .A2(\output_c[10][25] ),
    .A3(_1374_),
    .A4(_1375_),
    .B1(\output_c[10][27] ),
    .X(_1376_));
 sky130_fd_sc_hd__and2b_1 _2811_ (.A_N(_1371_),
    .B(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _2812_ (.A(_1377_),
    .X(_0933_));
 sky130_fd_sc_hd__and2_1 _2813_ (.A(_1358_),
    .B(_1365_),
    .X(_1378_));
 sky130_fd_sc_hd__and4_1 _2814_ (.A(\output_c[10][25] ),
    .B(_1374_),
    .C(_1355_),
    .D(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__xor2_1 _2815_ (.A(net109),
    .B(_1379_),
    .X(_0932_));
 sky130_fd_sc_hd__a21o_1 _2816_ (.A1(_1374_),
    .A2(_1375_),
    .B1(\output_c[10][25] ),
    .X(_1380_));
 sky130_fd_sc_hd__and2b_1 _2817_ (.A_N(_1379_),
    .B(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _2818_ (.A(_1381_),
    .X(_0931_));
 sky130_fd_sc_hd__xor2_1 _2819_ (.A(_1374_),
    .B(_1375_),
    .X(_0930_));
 sky130_fd_sc_hd__buf_1 _2820_ (.A(_1378_),
    .X(_1382_));
 sky130_fd_sc_hd__a31o_1 _2821_ (.A1(\output_c[10][22] ),
    .A2(_1353_),
    .A3(_1382_),
    .B1(net485),
    .X(_1383_));
 sky130_fd_sc_hd__a21boi_1 _2822_ (.A1(_1355_),
    .A2(_1382_),
    .B1_N(_1383_),
    .Y(_0929_));
 sky130_fd_sc_hd__and3_1 _2823_ (.A(_1352_),
    .B(_1359_),
    .C(_1370_),
    .X(_1384_));
 sky130_fd_sc_hd__and3_1 _2824_ (.A(\output_c[10][21] ),
    .B(\output_c[10][20] ),
    .C(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__xor2_1 _2825_ (.A(net181),
    .B(_1385_),
    .X(_0928_));
 sky130_fd_sc_hd__a21oi_1 _2826_ (.A1(net234),
    .A2(_1384_),
    .B1(net247),
    .Y(_1386_));
 sky130_fd_sc_hd__nor2_1 _2827_ (.A(_1385_),
    .B(_1386_),
    .Y(_0927_));
 sky130_fd_sc_hd__xor2_1 _2828_ (.A(net234),
    .B(_1384_),
    .X(_0926_));
 sky130_fd_sc_hd__and3_1 _2829_ (.A(\output_c[10][16] ),
    .B(_1359_),
    .C(_1370_),
    .X(_1387_));
 sky130_fd_sc_hd__a31o_1 _2830_ (.A1(\output_c[10][18] ),
    .A2(\output_c[10][17] ),
    .A3(_1387_),
    .B1(\output_c[10][19] ),
    .X(_1388_));
 sky130_fd_sc_hd__and2b_1 _2831_ (.A_N(_1384_),
    .B(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _2832_ (.A(_1389_),
    .X(_0925_));
 sky130_fd_sc_hd__and3_1 _2833_ (.A(\output_c[10][17] ),
    .B(\output_c[10][16] ),
    .C(_1382_),
    .X(_1390_));
 sky130_fd_sc_hd__xor2_1 _2834_ (.A(net182),
    .B(_1390_),
    .X(_0924_));
 sky130_fd_sc_hd__nor2_1 _2835_ (.A(net476),
    .B(_1387_),
    .Y(_1391_));
 sky130_fd_sc_hd__nor2_1 _2836_ (.A(_1390_),
    .B(_1391_),
    .Y(_0923_));
 sky130_fd_sc_hd__xor2_1 _2837_ (.A(net210),
    .B(_1382_),
    .X(_0922_));
 sky130_fd_sc_hd__and3_1 _2838_ (.A(\output_c[10][12] ),
    .B(_1356_),
    .C(_1365_),
    .X(_1392_));
 sky130_fd_sc_hd__and3_1 _2839_ (.A(\output_c[10][14] ),
    .B(\output_c[10][13] ),
    .C(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__xor2_1 _2840_ (.A(net51),
    .B(_1393_),
    .X(_0921_));
 sky130_fd_sc_hd__buf_1 _2841_ (.A(_1370_),
    .X(_1394_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2842_ (.A(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__a21oi_1 _2843_ (.A1(_1357_),
    .A2(_1395_),
    .B1(net206),
    .Y(_1396_));
 sky130_fd_sc_hd__nor2_1 _2844_ (.A(_1393_),
    .B(_1396_),
    .Y(_0920_));
 sky130_fd_sc_hd__nor2_1 _2845_ (.A(net354),
    .B(_1392_),
    .Y(_1397_));
 sky130_fd_sc_hd__a21oi_1 _2846_ (.A1(_1357_),
    .A2(_1395_),
    .B1(_1397_),
    .Y(_0919_));
 sky130_fd_sc_hd__and2_1 _2847_ (.A(_1356_),
    .B(_1394_),
    .X(_1398_));
 sky130_fd_sc_hd__nor2_1 _2848_ (.A(net295),
    .B(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__nor2_1 _2849_ (.A(_1392_),
    .B(_1399_),
    .Y(_0918_));
 sky130_fd_sc_hd__and3_1 _2850_ (.A(\output_c[10][9] ),
    .B(\output_c[10][8] ),
    .C(_1394_),
    .X(_1400_));
 sky130_fd_sc_hd__a21oi_1 _2851_ (.A1(\output_c[10][10] ),
    .A2(_1400_),
    .B1(net156),
    .Y(_1401_));
 sky130_fd_sc_hd__nor2_1 _2852_ (.A(_1398_),
    .B(net157),
    .Y(_0917_));
 sky130_fd_sc_hd__xor2_1 _2853_ (.A(net174),
    .B(_1400_),
    .X(_0916_));
 sky130_fd_sc_hd__a21oi_1 _2854_ (.A1(\output_c[10][8] ),
    .A2(_1395_),
    .B1(net204),
    .Y(_1402_));
 sky130_fd_sc_hd__nor2_1 _2855_ (.A(_1400_),
    .B(net205),
    .Y(_0915_));
 sky130_fd_sc_hd__xor2_1 _2856_ (.A(net252),
    .B(_1395_),
    .X(_0914_));
 sky130_fd_sc_hd__buf_1 _2857_ (.A(_1363_),
    .X(_1403_));
 sky130_fd_sc_hd__and3_1 _2858_ (.A(\output_c[10][5] ),
    .B(_1360_),
    .C(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__a21o_1 _2859_ (.A1(\output_c[10][6] ),
    .A2(_1404_),
    .B1(\output_c[10][7] ),
    .X(_1405_));
 sky130_fd_sc_hd__and2b_1 _2860_ (.A_N(_1394_),
    .B(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _2861_ (.A(_1406_),
    .X(_0913_));
 sky130_fd_sc_hd__xor2_1 _2862_ (.A(net358),
    .B(_1404_),
    .X(_0912_));
 sky130_fd_sc_hd__a21oi_1 _2863_ (.A1(_1360_),
    .A2(_1403_),
    .B1(net480),
    .Y(_1407_));
 sky130_fd_sc_hd__nor2_1 _2864_ (.A(_1404_),
    .B(_1407_),
    .Y(_0911_));
 sky130_fd_sc_hd__xor2_1 _2865_ (.A(_1360_),
    .B(_1403_),
    .X(_0910_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2866_ (.A(_1154_),
    .X(_1408_));
 sky130_fd_sc_hd__and3_1 _2867_ (.A(\output_c[10][1] ),
    .B(_1408_),
    .C(_1361_),
    .X(_1409_));
 sky130_fd_sc_hd__and2_1 _2868_ (.A(\output_c[10][2] ),
    .B(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__o21ba_1 _2869_ (.A1(net404),
    .A2(_1410_),
    .B1_N(_1403_),
    .X(_0909_));
 sky130_fd_sc_hd__nor2_1 _2870_ (.A(net462),
    .B(_1409_),
    .Y(_1411_));
 sky130_fd_sc_hd__nor2_1 _2871_ (.A(_1410_),
    .B(_1411_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21oi_1 _2872_ (.A1(_1346_),
    .A2(_1361_),
    .B1(net436),
    .Y(_1412_));
 sky130_fd_sc_hd__nor2_1 _2873_ (.A(_1409_),
    .B(_1412_),
    .Y(_0907_));
 sky130_fd_sc_hd__buf_1 _2874_ (.A(_1147_),
    .X(_1413_));
 sky130_fd_sc_hd__buf_1 _2875_ (.A(_1155_),
    .X(_1414_));
 sky130_fd_sc_hd__and3_1 _2876_ (.A(_1349_),
    .B(\input_a[10][0] ),
    .C(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__o2bb2a_1 _2877_ (.A1_N(_1413_),
    .A2_N(_1361_),
    .B1(_1415_),
    .B2(net168),
    .X(_0906_));
 sky130_fd_sc_hd__and4_1 _2878_ (.A(\output_c[9][27] ),
    .B(\output_c[9][26] ),
    .C(\output_c[9][25] ),
    .D(\output_c[9][24] ),
    .X(_1416_));
 sky130_fd_sc_hd__and4_1 _2879_ (.A(\output_c[9][19] ),
    .B(\output_c[9][18] ),
    .C(\output_c[9][17] ),
    .D(\output_c[9][16] ),
    .X(_1417_));
 sky130_fd_sc_hd__and3_1 _2880_ (.A(\output_c[9][21] ),
    .B(\output_c[9][20] ),
    .C(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__and3_1 _2881_ (.A(\output_c[9][23] ),
    .B(\output_c[9][22] ),
    .C(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__and4_1 _2882_ (.A(\output_c[9][11] ),
    .B(\output_c[9][10] ),
    .C(\output_c[9][9] ),
    .D(\output_c[9][8] ),
    .X(_1420_));
 sky130_fd_sc_hd__and3_1 _2883_ (.A(\output_c[9][13] ),
    .B(\output_c[9][12] ),
    .C(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__and3_1 _2884_ (.A(\output_c[9][15] ),
    .B(\output_c[9][14] ),
    .C(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__buf_1 _2885_ (.A(\output_c[9][4] ),
    .X(_1423_));
 sky130_fd_sc_hd__buf_1 _2886_ (.A(\input_b[15][0] ),
    .X(_1424_));
 sky130_fd_sc_hd__and3_1 _2887_ (.A(\output_c[9][0] ),
    .B(_1424_),
    .C(\input_a[9][0] ),
    .X(_1425_));
 sky130_fd_sc_hd__and2_1 _2888_ (.A(\output_c[9][3] ),
    .B(\output_c[9][2] ),
    .X(_1426_));
 sky130_fd_sc_hd__and4_1 _2889_ (.A(\output_c[9][1] ),
    .B(_1079_),
    .C(_1425_),
    .D(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__and2_1 _2890_ (.A(\output_c[9][7] ),
    .B(\output_c[9][6] ),
    .X(_1428_));
 sky130_fd_sc_hd__and4_1 _2891_ (.A(\output_c[9][5] ),
    .B(_1423_),
    .C(_1427_),
    .D(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__and4_1 _2892_ (.A(_1416_),
    .B(_1419_),
    .C(_1422_),
    .D(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__and4_1 _2893_ (.A(\output_c[9][30] ),
    .B(\output_c[9][29] ),
    .C(\output_c[9][28] ),
    .D(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__xor2_1 _2894_ (.A(net43),
    .B(_1431_),
    .X(_0905_));
 sky130_fd_sc_hd__and2_1 _2895_ (.A(\output_c[9][6] ),
    .B(\output_c[9][5] ),
    .X(_1432_));
 sky130_fd_sc_hd__and4_1 _2896_ (.A(\output_c[9][7] ),
    .B(\output_c[9][4] ),
    .C(_1427_),
    .D(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__and4_1 _2897_ (.A(_1416_),
    .B(_1419_),
    .C(_1422_),
    .D(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__and3_1 _2898_ (.A(\output_c[9][29] ),
    .B(\output_c[9][28] ),
    .C(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__xor2_1 _2899_ (.A(net76),
    .B(_1435_),
    .X(_0904_));
 sky130_fd_sc_hd__a21oi_1 _2900_ (.A1(net265),
    .A2(_1434_),
    .B1(net318),
    .Y(_1436_));
 sky130_fd_sc_hd__nor2_1 _2901_ (.A(_1435_),
    .B(_1436_),
    .Y(_0903_));
 sky130_fd_sc_hd__xor2_1 _2902_ (.A(net265),
    .B(_1434_),
    .X(_0902_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2903_ (.A(\output_c[9][24] ),
    .X(_1437_));
 sky130_fd_sc_hd__and3_1 _2904_ (.A(_1419_),
    .B(_1422_),
    .C(_1433_),
    .X(_1438_));
 sky130_fd_sc_hd__a41o_1 _2905_ (.A1(\output_c[9][26] ),
    .A2(\output_c[9][25] ),
    .A3(_1437_),
    .A4(_1438_),
    .B1(\output_c[9][27] ),
    .X(_1439_));
 sky130_fd_sc_hd__and2b_1 _2906_ (.A_N(_1434_),
    .B(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _2907_ (.A(_1440_),
    .X(_0901_));
 sky130_fd_sc_hd__buf_1 _2908_ (.A(_1438_),
    .X(_1441_));
 sky130_fd_sc_hd__nand3_1 _2909_ (.A(\output_c[9][25] ),
    .B(_1437_),
    .C(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__xnor2_1 _2910_ (.A(net137),
    .B(_1442_),
    .Y(_0900_));
 sky130_fd_sc_hd__a21o_1 _2911_ (.A1(_1437_),
    .A2(_1441_),
    .B1(\output_c[9][25] ),
    .X(_1443_));
 sky130_fd_sc_hd__and2_1 _2912_ (.A(_1442_),
    .B(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _2913_ (.A(_1444_),
    .X(_0899_));
 sky130_fd_sc_hd__xor2_1 _2914_ (.A(_1437_),
    .B(_1441_),
    .X(_0898_));
 sky130_fd_sc_hd__buf_1 _2915_ (.A(_1422_),
    .X(_1445_));
 sky130_fd_sc_hd__a41o_1 _2916_ (.A1(\output_c[9][22] ),
    .A2(_1418_),
    .A3(_1445_),
    .A4(_1429_),
    .B1(\output_c[9][23] ),
    .X(_1446_));
 sky130_fd_sc_hd__and2b_1 _2917_ (.A_N(_1441_),
    .B(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _2918_ (.A(_1447_),
    .X(_0897_));
 sky130_fd_sc_hd__buf_1 _2919_ (.A(_1433_),
    .X(_1448_));
 sky130_fd_sc_hd__and3_1 _2920_ (.A(_1417_),
    .B(_1445_),
    .C(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__and3_1 _2921_ (.A(\output_c[9][21] ),
    .B(\output_c[9][20] ),
    .C(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__xor2_1 _2922_ (.A(net110),
    .B(_1450_),
    .X(_0896_));
 sky130_fd_sc_hd__a21oi_1 _2923_ (.A1(net280),
    .A2(_1449_),
    .B1(net346),
    .Y(_1451_));
 sky130_fd_sc_hd__nor2_1 _2924_ (.A(_1450_),
    .B(_1451_),
    .Y(_0895_));
 sky130_fd_sc_hd__xor2_1 _2925_ (.A(net280),
    .B(_1449_),
    .X(_0894_));
 sky130_fd_sc_hd__and3_1 _2926_ (.A(\output_c[9][16] ),
    .B(_1445_),
    .C(_1448_),
    .X(_1452_));
 sky130_fd_sc_hd__and3_1 _2927_ (.A(\output_c[9][18] ),
    .B(\output_c[9][17] ),
    .C(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__o21ba_1 _2928_ (.A1(net147),
    .A2(_1453_),
    .B1_N(_1449_),
    .X(_0893_));
 sky130_fd_sc_hd__a21oi_1 _2929_ (.A1(net246),
    .A2(_1452_),
    .B1(net306),
    .Y(_1454_));
 sky130_fd_sc_hd__nor2_1 _2930_ (.A(_1453_),
    .B(_1454_),
    .Y(_0892_));
 sky130_fd_sc_hd__xor2_1 _2931_ (.A(net246),
    .B(_1452_),
    .X(_0891_));
 sky130_fd_sc_hd__buf_1 _2932_ (.A(_1448_),
    .X(_1455_));
 sky130_fd_sc_hd__a21o_1 _2933_ (.A1(_1445_),
    .A2(_1455_),
    .B1(\output_c[9][16] ),
    .X(_1456_));
 sky130_fd_sc_hd__and2b_1 _2934_ (.A_N(_1452_),
    .B(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _2935_ (.A(_1457_),
    .X(_0890_));
 sky130_fd_sc_hd__and3_1 _2936_ (.A(\output_c[9][12] ),
    .B(_1420_),
    .C(_1429_),
    .X(_1458_));
 sky130_fd_sc_hd__and3_1 _2937_ (.A(\output_c[9][14] ),
    .B(\output_c[9][13] ),
    .C(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__xor2_1 _2938_ (.A(net54),
    .B(_1459_),
    .X(_0889_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2939_ (.A(_1455_),
    .X(_1460_));
 sky130_fd_sc_hd__a21oi_1 _2940_ (.A1(_1421_),
    .A2(_1460_),
    .B1(net238),
    .Y(_1461_));
 sky130_fd_sc_hd__nor2_1 _2941_ (.A(_1459_),
    .B(_1461_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor2_1 _2942_ (.A(net230),
    .B(_1458_),
    .Y(_1462_));
 sky130_fd_sc_hd__a21oi_1 _2943_ (.A1(_1421_),
    .A2(_1460_),
    .B1(_1462_),
    .Y(_0887_));
 sky130_fd_sc_hd__and2_1 _2944_ (.A(_1420_),
    .B(_1455_),
    .X(_1463_));
 sky130_fd_sc_hd__nor2_1 _2945_ (.A(net325),
    .B(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__nor2_1 _2946_ (.A(_1458_),
    .B(_1464_),
    .Y(_0886_));
 sky130_fd_sc_hd__and3_1 _2947_ (.A(\output_c[9][9] ),
    .B(\output_c[9][8] ),
    .C(_1448_),
    .X(_1465_));
 sky130_fd_sc_hd__a21oi_1 _2948_ (.A1(\output_c[9][10] ),
    .A2(_1465_),
    .B1(net94),
    .Y(_1466_));
 sky130_fd_sc_hd__nor2_1 _2949_ (.A(_1463_),
    .B(net95),
    .Y(_0885_));
 sky130_fd_sc_hd__xor2_1 _2950_ (.A(net128),
    .B(_1465_),
    .X(_0884_));
 sky130_fd_sc_hd__a21oi_1 _2951_ (.A1(\output_c[9][8] ),
    .A2(_1460_),
    .B1(net290),
    .Y(_1467_));
 sky130_fd_sc_hd__nor2_1 _2952_ (.A(_1465_),
    .B(net291),
    .Y(_0883_));
 sky130_fd_sc_hd__xor2_1 _2953_ (.A(net305),
    .B(_1460_),
    .X(_0882_));
 sky130_fd_sc_hd__buf_1 _2954_ (.A(_1427_),
    .X(_1468_));
 sky130_fd_sc_hd__and3_1 _2955_ (.A(\output_c[9][5] ),
    .B(_1423_),
    .C(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__a21o_1 _2956_ (.A1(\output_c[9][6] ),
    .A2(_1469_),
    .B1(\output_c[9][7] ),
    .X(_1470_));
 sky130_fd_sc_hd__and2b_1 _2957_ (.A_N(_1455_),
    .B(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _2958_ (.A(_1471_),
    .X(_0881_));
 sky130_fd_sc_hd__xor2_1 _2959_ (.A(net276),
    .B(_1469_),
    .X(_0880_));
 sky130_fd_sc_hd__a21oi_1 _2960_ (.A1(_1423_),
    .A2(_1468_),
    .B1(net455),
    .Y(_1472_));
 sky130_fd_sc_hd__nor2_1 _2961_ (.A(_1469_),
    .B(_1472_),
    .Y(_0879_));
 sky130_fd_sc_hd__xor2_1 _2962_ (.A(_1423_),
    .B(_1468_),
    .X(_0878_));
 sky130_fd_sc_hd__and3_1 _2963_ (.A(\output_c[9][1] ),
    .B(_1408_),
    .C(_1425_),
    .X(_1473_));
 sky130_fd_sc_hd__and2_1 _2964_ (.A(\output_c[9][2] ),
    .B(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__o21ba_1 _2965_ (.A1(net197),
    .A2(_1474_),
    .B1_N(_1468_),
    .X(_0877_));
 sky130_fd_sc_hd__nor2_1 _2966_ (.A(net446),
    .B(_1473_),
    .Y(_1475_));
 sky130_fd_sc_hd__nor2_1 _2967_ (.A(_1474_),
    .B(_1475_),
    .Y(_0876_));
 sky130_fd_sc_hd__a21oi_1 _2968_ (.A1(_1346_),
    .A2(_1425_),
    .B1(net330),
    .Y(_1476_));
 sky130_fd_sc_hd__nor2_1 _2969_ (.A(_1473_),
    .B(_1476_),
    .Y(_0875_));
 sky130_fd_sc_hd__and3_1 _2970_ (.A(_1349_),
    .B(\input_a[9][0] ),
    .C(_1414_),
    .X(_1477_));
 sky130_fd_sc_hd__o2bb2a_1 _2971_ (.A1_N(_1413_),
    .A2_N(_1425_),
    .B1(_1477_),
    .B2(net155),
    .X(_0874_));
 sky130_fd_sc_hd__and2_1 _2972_ (.A(\output_c[8][25] ),
    .B(\output_c[8][24] ),
    .X(_1478_));
 sky130_fd_sc_hd__and3_1 _2973_ (.A(\output_c[8][27] ),
    .B(\output_c[8][26] ),
    .C(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__and4_1 _2974_ (.A(\output_c[8][19] ),
    .B(\output_c[8][18] ),
    .C(\output_c[8][17] ),
    .D(\output_c[8][16] ),
    .X(_1480_));
 sky130_fd_sc_hd__and3_1 _2975_ (.A(\output_c[8][21] ),
    .B(\output_c[8][20] ),
    .C(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__and3_1 _2976_ (.A(\output_c[8][23] ),
    .B(\output_c[8][22] ),
    .C(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__and4_1 _2977_ (.A(\output_c[8][11] ),
    .B(\output_c[8][10] ),
    .C(\output_c[8][9] ),
    .D(\output_c[8][8] ),
    .X(_1483_));
 sky130_fd_sc_hd__and3_1 _2978_ (.A(\output_c[8][15] ),
    .B(\output_c[8][14] ),
    .C(\output_c[8][13] ),
    .X(_1484_));
 sky130_fd_sc_hd__and3_1 _2979_ (.A(\output_c[8][12] ),
    .B(_1483_),
    .C(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__buf_1 _2980_ (.A(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__buf_1 _2981_ (.A(\input_b[15][0] ),
    .X(_1487_));
 sky130_fd_sc_hd__and3_1 _2982_ (.A(\output_c[8][0] ),
    .B(_1487_),
    .C(\input_a[8][0] ),
    .X(_1488_));
 sky130_fd_sc_hd__and2_1 _2983_ (.A(\output_c[8][3] ),
    .B(\output_c[8][2] ),
    .X(_1489_));
 sky130_fd_sc_hd__and4_1 _2984_ (.A(\output_c[8][1] ),
    .B(_1101_),
    .C(_1488_),
    .D(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__and2_1 _2985_ (.A(\output_c[8][7] ),
    .B(\output_c[8][6] ),
    .X(_1491_));
 sky130_fd_sc_hd__and4_1 _2986_ (.A(\output_c[8][5] ),
    .B(\output_c[8][4] ),
    .C(_1490_),
    .D(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__and4_1 _2987_ (.A(_1479_),
    .B(_1482_),
    .C(_1486_),
    .D(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__and4_1 _2988_ (.A(\output_c[8][30] ),
    .B(\output_c[8][29] ),
    .C(\output_c[8][28] ),
    .D(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__xor2_1 _2989_ (.A(net40),
    .B(_1494_),
    .X(_0873_));
 sky130_fd_sc_hd__buf_1 _2990_ (.A(\output_c[8][4] ),
    .X(_1495_));
 sky130_fd_sc_hd__and2_1 _2991_ (.A(\output_c[8][6] ),
    .B(\output_c[8][5] ),
    .X(_1496_));
 sky130_fd_sc_hd__and4_1 _2992_ (.A(\output_c[8][7] ),
    .B(_1495_),
    .C(_1490_),
    .D(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__and4_2 _2993_ (.A(_1479_),
    .B(_1482_),
    .C(_1485_),
    .D(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__and3_1 _2994_ (.A(\output_c[8][29] ),
    .B(\output_c[8][28] ),
    .C(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__xor2_1 _2995_ (.A(net82),
    .B(_1499_),
    .X(_0872_));
 sky130_fd_sc_hd__a21oi_1 _2996_ (.A1(net273),
    .A2(_1498_),
    .B1(net333),
    .Y(_1500_));
 sky130_fd_sc_hd__nor2_1 _2997_ (.A(_1499_),
    .B(_1500_),
    .Y(_0871_));
 sky130_fd_sc_hd__xor2_1 _2998_ (.A(net273),
    .B(_1498_),
    .X(_0870_));
 sky130_fd_sc_hd__buf_1 _2999_ (.A(_1482_),
    .X(_1501_));
 sky130_fd_sc_hd__buf_1 _3000_ (.A(_1497_),
    .X(_1502_));
 sky130_fd_sc_hd__and4_1 _3001_ (.A(_1478_),
    .B(_1501_),
    .C(_1486_),
    .D(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__a21oi_1 _3002_ (.A1(\output_c[8][26] ),
    .A2(_1503_),
    .B1(net202),
    .Y(_1504_));
 sky130_fd_sc_hd__nor2_1 _3003_ (.A(_1498_),
    .B(net203),
    .Y(_0869_));
 sky130_fd_sc_hd__xor2_1 _3004_ (.A(net259),
    .B(_1503_),
    .X(_0868_));
 sky130_fd_sc_hd__and2_1 _3005_ (.A(_1485_),
    .B(_1492_),
    .X(_1505_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3006_ (.A(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__nand3_1 _3007_ (.A(\output_c[8][24] ),
    .B(_1501_),
    .C(_1506_),
    .Y(_1507_));
 sky130_fd_sc_hd__xnor2_1 _3008_ (.A(net78),
    .B(_1507_),
    .Y(_0867_));
 sky130_fd_sc_hd__a31o_1 _3009_ (.A1(_1501_),
    .A2(_1486_),
    .A3(_1502_),
    .B1(\output_c[8][24] ),
    .X(_1508_));
 sky130_fd_sc_hd__and2_1 _3010_ (.A(_1507_),
    .B(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _3011_ (.A(_1509_),
    .X(_0866_));
 sky130_fd_sc_hd__a31o_1 _3012_ (.A1(\output_c[8][22] ),
    .A2(_1481_),
    .A3(_1506_),
    .B1(net484),
    .X(_1510_));
 sky130_fd_sc_hd__a21boi_1 _3013_ (.A1(_1501_),
    .A2(_1506_),
    .B1_N(_1510_),
    .Y(_0865_));
 sky130_fd_sc_hd__and3_1 _3014_ (.A(_1480_),
    .B(_1486_),
    .C(_1497_),
    .X(_1511_));
 sky130_fd_sc_hd__and3_1 _3015_ (.A(\output_c[8][21] ),
    .B(\output_c[8][20] ),
    .C(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__xor2_1 _3016_ (.A(net220),
    .B(_1512_),
    .X(_0864_));
 sky130_fd_sc_hd__a21oi_1 _3017_ (.A1(net415),
    .A2(_1511_),
    .B1(net437),
    .Y(_1513_));
 sky130_fd_sc_hd__nor2_1 _3018_ (.A(_1512_),
    .B(_1513_),
    .Y(_0863_));
 sky130_fd_sc_hd__xor2_1 _3019_ (.A(net415),
    .B(_1511_),
    .X(_0862_));
 sky130_fd_sc_hd__and3_1 _3020_ (.A(\output_c[8][16] ),
    .B(_1485_),
    .C(_1497_),
    .X(_1514_));
 sky130_fd_sc_hd__a31o_1 _3021_ (.A1(\output_c[8][18] ),
    .A2(\output_c[8][17] ),
    .A3(_1514_),
    .B1(\output_c[8][19] ),
    .X(_1515_));
 sky130_fd_sc_hd__and2b_1 _3022_ (.A_N(_1511_),
    .B(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3023_ (.A(_1516_),
    .X(_0861_));
 sky130_fd_sc_hd__and3_1 _3024_ (.A(\output_c[8][17] ),
    .B(\output_c[8][16] ),
    .C(_1505_),
    .X(_1517_));
 sky130_fd_sc_hd__xor2_1 _3025_ (.A(net199),
    .B(_1517_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _3026_ (.A(net469),
    .B(_1514_),
    .Y(_1518_));
 sky130_fd_sc_hd__nor2_1 _3027_ (.A(_1517_),
    .B(_1518_),
    .Y(_0859_));
 sky130_fd_sc_hd__xor2_1 _3028_ (.A(net185),
    .B(_1506_),
    .X(_0858_));
 sky130_fd_sc_hd__and3_1 _3029_ (.A(\output_c[8][12] ),
    .B(_1483_),
    .C(_1492_),
    .X(_1519_));
 sky130_fd_sc_hd__and3_1 _3030_ (.A(\output_c[8][14] ),
    .B(\output_c[8][13] ),
    .C(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__xor2_1 _3031_ (.A(net56),
    .B(_1520_),
    .X(_0857_));
 sky130_fd_sc_hd__a21o_1 _3032_ (.A1(\output_c[8][13] ),
    .A2(_1519_),
    .B1(\output_c[8][14] ),
    .X(_1521_));
 sky130_fd_sc_hd__and2b_1 _3033_ (.A_N(_1520_),
    .B(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3034_ (.A(_1522_),
    .X(_0856_));
 sky130_fd_sc_hd__xor2_1 _3035_ (.A(net431),
    .B(_1519_),
    .X(_0855_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3036_ (.A(_1502_),
    .X(_1523_));
 sky130_fd_sc_hd__and2_1 _3037_ (.A(_1483_),
    .B(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__nor2_1 _3038_ (.A(net360),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nor2_1 _3039_ (.A(_1519_),
    .B(_1525_),
    .Y(_0854_));
 sky130_fd_sc_hd__and3_1 _3040_ (.A(\output_c[8][9] ),
    .B(\output_c[8][8] ),
    .C(_1502_),
    .X(_1526_));
 sky130_fd_sc_hd__a21oi_1 _3041_ (.A1(net105),
    .A2(_1526_),
    .B1(net141),
    .Y(_1527_));
 sky130_fd_sc_hd__nor2_1 _3042_ (.A(_1524_),
    .B(_1527_),
    .Y(_0853_));
 sky130_fd_sc_hd__xor2_1 _3043_ (.A(net105),
    .B(_1526_),
    .X(_0852_));
 sky130_fd_sc_hd__a21oi_1 _3044_ (.A1(\output_c[8][8] ),
    .A2(_1523_),
    .B1(net253),
    .Y(_1528_));
 sky130_fd_sc_hd__nor2_1 _3045_ (.A(_1526_),
    .B(net254),
    .Y(_0851_));
 sky130_fd_sc_hd__xor2_1 _3046_ (.A(net270),
    .B(_1523_),
    .X(_0850_));
 sky130_fd_sc_hd__buf_1 _3047_ (.A(_1490_),
    .X(_1529_));
 sky130_fd_sc_hd__and3_1 _3048_ (.A(\output_c[8][5] ),
    .B(_1495_),
    .C(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__a21o_1 _3049_ (.A1(\output_c[8][6] ),
    .A2(_1530_),
    .B1(\output_c[8][7] ),
    .X(_1531_));
 sky130_fd_sc_hd__and2b_1 _3050_ (.A_N(_1523_),
    .B(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3051_ (.A(_1532_),
    .X(_0849_));
 sky130_fd_sc_hd__xor2_1 _3052_ (.A(net287),
    .B(_1530_),
    .X(_0848_));
 sky130_fd_sc_hd__a21oi_1 _3053_ (.A1(_1495_),
    .A2(_1529_),
    .B1(net466),
    .Y(_1533_));
 sky130_fd_sc_hd__nor2_1 _3054_ (.A(_1530_),
    .B(_1533_),
    .Y(_0847_));
 sky130_fd_sc_hd__xor2_1 _3055_ (.A(_1495_),
    .B(_1529_),
    .X(_0846_));
 sky130_fd_sc_hd__and3_1 _3056_ (.A(\output_c[8][1] ),
    .B(_1408_),
    .C(_1488_),
    .X(_1534_));
 sky130_fd_sc_hd__and2_1 _3057_ (.A(\output_c[8][2] ),
    .B(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__o21ba_1 _3058_ (.A1(net218),
    .A2(_1535_),
    .B1_N(_1529_),
    .X(_0845_));
 sky130_fd_sc_hd__nor2_1 _3059_ (.A(net428),
    .B(_1534_),
    .Y(_1536_));
 sky130_fd_sc_hd__nor2_1 _3060_ (.A(_1535_),
    .B(_1536_),
    .Y(_0844_));
 sky130_fd_sc_hd__a21oi_1 _3061_ (.A1(_1346_),
    .A2(_1488_),
    .B1(net384),
    .Y(_1537_));
 sky130_fd_sc_hd__nor2_1 _3062_ (.A(_1534_),
    .B(_1537_),
    .Y(_0843_));
 sky130_fd_sc_hd__and3_1 _3063_ (.A(_1349_),
    .B(\input_a[8][0] ),
    .C(_1414_),
    .X(_1538_));
 sky130_fd_sc_hd__o2bb2a_1 _3064_ (.A1_N(_1413_),
    .A2_N(_1488_),
    .B1(_1538_),
    .B2(net208),
    .X(_0842_));
 sky130_fd_sc_hd__and2_1 _3065_ (.A(\output_c[7][25] ),
    .B(\output_c[7][24] ),
    .X(_1539_));
 sky130_fd_sc_hd__and3_1 _3066_ (.A(\output_c[7][27] ),
    .B(\output_c[7][26] ),
    .C(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__and4_1 _3067_ (.A(\output_c[7][19] ),
    .B(\output_c[7][18] ),
    .C(\output_c[7][17] ),
    .D(\output_c[7][16] ),
    .X(_1541_));
 sky130_fd_sc_hd__and3_1 _3068_ (.A(\output_c[7][21] ),
    .B(\output_c[7][20] ),
    .C(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__and3_1 _3069_ (.A(\output_c[7][23] ),
    .B(\output_c[7][22] ),
    .C(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__and4_1 _3070_ (.A(\output_c[7][11] ),
    .B(\output_c[7][10] ),
    .C(\output_c[7][9] ),
    .D(\output_c[7][8] ),
    .X(_1544_));
 sky130_fd_sc_hd__and3_1 _3071_ (.A(\output_c[7][15] ),
    .B(\output_c[7][14] ),
    .C(\output_c[7][13] ),
    .X(_1545_));
 sky130_fd_sc_hd__and3_1 _3072_ (.A(\output_c[7][12] ),
    .B(_1544_),
    .C(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__buf_1 _3073_ (.A(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__and3_1 _3074_ (.A(\output_c[7][0] ),
    .B(_1487_),
    .C(\input_a[7][0] ),
    .X(_1548_));
 sky130_fd_sc_hd__and2_1 _3075_ (.A(\output_c[7][3] ),
    .B(\output_c[7][2] ),
    .X(_1549_));
 sky130_fd_sc_hd__and4_1 _3076_ (.A(\output_c[7][1] ),
    .B(_1101_),
    .C(_1548_),
    .D(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__and2_1 _3077_ (.A(\output_c[7][7] ),
    .B(\output_c[7][6] ),
    .X(_1551_));
 sky130_fd_sc_hd__and4_1 _3078_ (.A(\output_c[7][5] ),
    .B(\output_c[7][4] ),
    .C(_1550_),
    .D(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__and4_1 _3079_ (.A(_1540_),
    .B(_1543_),
    .C(_1547_),
    .D(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__and4_1 _3080_ (.A(\output_c[7][30] ),
    .B(\output_c[7][29] ),
    .C(\output_c[7][28] ),
    .D(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__xor2_1 _3081_ (.A(net49),
    .B(_1554_),
    .X(_0841_));
 sky130_fd_sc_hd__buf_1 _3082_ (.A(\output_c[7][4] ),
    .X(_1555_));
 sky130_fd_sc_hd__and2_1 _3083_ (.A(\output_c[7][6] ),
    .B(\output_c[7][5] ),
    .X(_1556_));
 sky130_fd_sc_hd__and4_1 _3084_ (.A(\output_c[7][7] ),
    .B(_1555_),
    .C(_1550_),
    .D(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__and4_1 _3085_ (.A(_1540_),
    .B(_1543_),
    .C(_1546_),
    .D(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__and3_1 _3086_ (.A(\output_c[7][29] ),
    .B(\output_c[7][28] ),
    .C(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__xor2_1 _3087_ (.A(net83),
    .B(_1559_),
    .X(_0840_));
 sky130_fd_sc_hd__a21oi_1 _3088_ (.A1(net399),
    .A2(_1558_),
    .B1(net432),
    .Y(_1560_));
 sky130_fd_sc_hd__nor2_1 _3089_ (.A(_1559_),
    .B(_1560_),
    .Y(_0839_));
 sky130_fd_sc_hd__xor2_1 _3090_ (.A(net399),
    .B(_1558_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_1 _3091_ (.A(_1543_),
    .X(_1561_));
 sky130_fd_sc_hd__buf_1 _3092_ (.A(_1557_),
    .X(_1562_));
 sky130_fd_sc_hd__and4_1 _3093_ (.A(_1539_),
    .B(_1561_),
    .C(_1547_),
    .D(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a21oi_1 _3094_ (.A1(net140),
    .A2(_1563_),
    .B1(net211),
    .Y(_1564_));
 sky130_fd_sc_hd__nor2_1 _3095_ (.A(_1558_),
    .B(_1564_),
    .Y(_0837_));
 sky130_fd_sc_hd__xor2_1 _3096_ (.A(net140),
    .B(_1563_),
    .X(_0836_));
 sky130_fd_sc_hd__and2_1 _3097_ (.A(_1546_),
    .B(_1552_),
    .X(_1565_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3098_ (.A(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__nand3_1 _3099_ (.A(\output_c[7][24] ),
    .B(_1561_),
    .C(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__xnor2_1 _3100_ (.A(net69),
    .B(_1567_),
    .Y(_0835_));
 sky130_fd_sc_hd__a31o_1 _3101_ (.A1(_1561_),
    .A2(_1547_),
    .A3(_1562_),
    .B1(\output_c[7][24] ),
    .X(_1568_));
 sky130_fd_sc_hd__and2_1 _3102_ (.A(_1567_),
    .B(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3103_ (.A(_1569_),
    .X(_0834_));
 sky130_fd_sc_hd__a31o_1 _3104_ (.A1(\output_c[7][22] ),
    .A2(_1542_),
    .A3(_1566_),
    .B1(net488),
    .X(_1570_));
 sky130_fd_sc_hd__a21boi_1 _3105_ (.A1(_1561_),
    .A2(_1566_),
    .B1_N(_1570_),
    .Y(_0833_));
 sky130_fd_sc_hd__and3_1 _3106_ (.A(_1541_),
    .B(_1547_),
    .C(_1557_),
    .X(_1571_));
 sky130_fd_sc_hd__and3_1 _3107_ (.A(\output_c[7][21] ),
    .B(\output_c[7][20] ),
    .C(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__xor2_1 _3108_ (.A(net151),
    .B(_1572_),
    .X(_0832_));
 sky130_fd_sc_hd__a21oi_1 _3109_ (.A1(net337),
    .A2(_1571_),
    .B1(net352),
    .Y(_1573_));
 sky130_fd_sc_hd__nor2_1 _3110_ (.A(_1572_),
    .B(_1573_),
    .Y(_0831_));
 sky130_fd_sc_hd__xor2_1 _3111_ (.A(net337),
    .B(_1571_),
    .X(_0830_));
 sky130_fd_sc_hd__and3_1 _3112_ (.A(\output_c[7][16] ),
    .B(_1546_),
    .C(_1557_),
    .X(_1574_));
 sky130_fd_sc_hd__a31o_1 _3113_ (.A1(\output_c[7][18] ),
    .A2(\output_c[7][17] ),
    .A3(_1574_),
    .B1(\output_c[7][19] ),
    .X(_1575_));
 sky130_fd_sc_hd__and2b_1 _3114_ (.A_N(_1571_),
    .B(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3115_ (.A(_1576_),
    .X(_0829_));
 sky130_fd_sc_hd__and3_1 _3116_ (.A(\output_c[7][17] ),
    .B(\output_c[7][16] ),
    .C(_1565_),
    .X(_1577_));
 sky130_fd_sc_hd__xor2_1 _3117_ (.A(net148),
    .B(_1577_),
    .X(_0828_));
 sky130_fd_sc_hd__nor2_1 _3118_ (.A(net483),
    .B(_1574_),
    .Y(_1578_));
 sky130_fd_sc_hd__nor2_1 _3119_ (.A(_1577_),
    .B(_1578_),
    .Y(_0827_));
 sky130_fd_sc_hd__xor2_1 _3120_ (.A(net241),
    .B(_1566_),
    .X(_0826_));
 sky130_fd_sc_hd__and3_1 _3121_ (.A(\output_c[7][12] ),
    .B(_1544_),
    .C(_1552_),
    .X(_1579_));
 sky130_fd_sc_hd__and3_1 _3122_ (.A(\output_c[7][14] ),
    .B(\output_c[7][13] ),
    .C(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__xor2_1 _3123_ (.A(net68),
    .B(_1580_),
    .X(_0825_));
 sky130_fd_sc_hd__a21o_1 _3124_ (.A1(\output_c[7][13] ),
    .A2(_1579_),
    .B1(\output_c[7][14] ),
    .X(_1581_));
 sky130_fd_sc_hd__and2b_1 _3125_ (.A_N(_1580_),
    .B(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _3126_ (.A(_1582_),
    .X(_0824_));
 sky130_fd_sc_hd__xor2_1 _3127_ (.A(net271),
    .B(_1579_),
    .X(_0823_));
 sky130_fd_sc_hd__buf_1 _3128_ (.A(_1562_),
    .X(_1583_));
 sky130_fd_sc_hd__and2_1 _3129_ (.A(_1544_),
    .B(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__nor2_1 _3130_ (.A(net292),
    .B(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__nor2_1 _3131_ (.A(_1579_),
    .B(_1585_),
    .Y(_0822_));
 sky130_fd_sc_hd__and3_1 _3132_ (.A(\output_c[7][9] ),
    .B(\output_c[7][8] ),
    .C(_1562_),
    .X(_1586_));
 sky130_fd_sc_hd__a21oi_1 _3133_ (.A1(\output_c[7][10] ),
    .A2(_1586_),
    .B1(net107),
    .Y(_1587_));
 sky130_fd_sc_hd__nor2_1 _3134_ (.A(_1584_),
    .B(net108),
    .Y(_0821_));
 sky130_fd_sc_hd__xor2_1 _3135_ (.A(net161),
    .B(_1586_),
    .X(_0820_));
 sky130_fd_sc_hd__a21oi_1 _3136_ (.A1(\output_c[7][8] ),
    .A2(_1583_),
    .B1(net281),
    .Y(_1588_));
 sky130_fd_sc_hd__nor2_1 _3137_ (.A(_1586_),
    .B(net282),
    .Y(_0819_));
 sky130_fd_sc_hd__xor2_1 _3138_ (.A(net364),
    .B(_1583_),
    .X(_0818_));
 sky130_fd_sc_hd__buf_1 _3139_ (.A(_1550_),
    .X(_1589_));
 sky130_fd_sc_hd__and3_1 _3140_ (.A(\output_c[7][5] ),
    .B(_1555_),
    .C(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__a21o_1 _3141_ (.A1(\output_c[7][6] ),
    .A2(_1590_),
    .B1(\output_c[7][7] ),
    .X(_1591_));
 sky130_fd_sc_hd__and2b_1 _3142_ (.A_N(_1583_),
    .B(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _3143_ (.A(_1592_),
    .X(_0817_));
 sky130_fd_sc_hd__xor2_1 _3144_ (.A(net300),
    .B(_1590_),
    .X(_0816_));
 sky130_fd_sc_hd__a21oi_1 _3145_ (.A1(_1555_),
    .A2(_1589_),
    .B1(net453),
    .Y(_1593_));
 sky130_fd_sc_hd__nor2_1 _3146_ (.A(_1590_),
    .B(_1593_),
    .Y(_0815_));
 sky130_fd_sc_hd__xor2_1 _3147_ (.A(_1555_),
    .B(_1589_),
    .X(_0814_));
 sky130_fd_sc_hd__and3_1 _3148_ (.A(\output_c[7][1] ),
    .B(_1408_),
    .C(_1548_),
    .X(_1594_));
 sky130_fd_sc_hd__and2_1 _3149_ (.A(\output_c[7][2] ),
    .B(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__o21ba_1 _3150_ (.A1(net249),
    .A2(_1595_),
    .B1_N(_1589_),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_1 _3151_ (.A(net472),
    .B(_1594_),
    .Y(_1596_));
 sky130_fd_sc_hd__nor2_1 _3152_ (.A(_1595_),
    .B(_1596_),
    .Y(_0812_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3153_ (.A(_1345_),
    .X(_1597_));
 sky130_fd_sc_hd__a21oi_1 _3154_ (.A1(_1597_),
    .A2(_1548_),
    .B1(net406),
    .Y(_1598_));
 sky130_fd_sc_hd__nor2_1 _3155_ (.A(_1594_),
    .B(_1598_),
    .Y(_0811_));
 sky130_fd_sc_hd__buf_1 _3156_ (.A(_1348_),
    .X(_1599_));
 sky130_fd_sc_hd__and3_1 _3157_ (.A(_1599_),
    .B(\input_a[7][0] ),
    .C(_1414_),
    .X(_1600_));
 sky130_fd_sc_hd__o2bb2a_1 _3158_ (.A1_N(_1413_),
    .A2_N(_1548_),
    .B1(_1600_),
    .B2(net216),
    .X(_0810_));
 sky130_fd_sc_hd__and4_1 _3159_ (.A(\output_c[6][27] ),
    .B(\output_c[6][26] ),
    .C(\output_c[6][25] ),
    .D(\output_c[6][24] ),
    .X(_1601_));
 sky130_fd_sc_hd__and4_1 _3160_ (.A(\output_c[6][19] ),
    .B(\output_c[6][18] ),
    .C(\output_c[6][17] ),
    .D(\output_c[6][16] ),
    .X(_1602_));
 sky130_fd_sc_hd__and3_1 _3161_ (.A(\output_c[6][21] ),
    .B(\output_c[6][20] ),
    .C(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__and3_1 _3162_ (.A(\output_c[6][23] ),
    .B(\output_c[6][22] ),
    .C(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__and4_1 _3163_ (.A(\output_c[6][11] ),
    .B(\output_c[6][10] ),
    .C(\output_c[6][9] ),
    .D(\output_c[6][8] ),
    .X(_1605_));
 sky130_fd_sc_hd__and3_1 _3164_ (.A(\output_c[6][13] ),
    .B(\output_c[6][12] ),
    .C(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__and3_1 _3165_ (.A(\output_c[6][15] ),
    .B(\output_c[6][14] ),
    .C(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__buf_1 _3166_ (.A(\output_c[6][4] ),
    .X(_1608_));
 sky130_fd_sc_hd__and3_1 _3167_ (.A(\output_c[6][0] ),
    .B(_1424_),
    .C(\input_a[6][0] ),
    .X(_1609_));
 sky130_fd_sc_hd__and2_1 _3168_ (.A(\output_c[6][3] ),
    .B(\output_c[6][2] ),
    .X(_1610_));
 sky130_fd_sc_hd__and4_1 _3169_ (.A(\output_c[6][1] ),
    .B(_1079_),
    .C(_1609_),
    .D(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__and2_1 _3170_ (.A(\output_c[6][7] ),
    .B(\output_c[6][6] ),
    .X(_1612_));
 sky130_fd_sc_hd__and4_1 _3171_ (.A(\output_c[6][5] ),
    .B(_1608_),
    .C(_1611_),
    .D(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__and4_1 _3172_ (.A(_1601_),
    .B(_1604_),
    .C(_1607_),
    .D(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__and4_1 _3173_ (.A(\output_c[6][30] ),
    .B(\output_c[6][29] ),
    .C(\output_c[6][28] ),
    .D(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__xor2_1 _3174_ (.A(net35),
    .B(_1615_),
    .X(_0809_));
 sky130_fd_sc_hd__and2_1 _3175_ (.A(\output_c[6][6] ),
    .B(\output_c[6][5] ),
    .X(_1616_));
 sky130_fd_sc_hd__and4_1 _3176_ (.A(\output_c[6][7] ),
    .B(\output_c[6][4] ),
    .C(_1611_),
    .D(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__and4_1 _3177_ (.A(_1601_),
    .B(_1604_),
    .C(_1607_),
    .D(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__and3_1 _3178_ (.A(\output_c[6][29] ),
    .B(\output_c[6][28] ),
    .C(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__xor2_1 _3179_ (.A(net75),
    .B(_1619_),
    .X(_0808_));
 sky130_fd_sc_hd__a21oi_1 _3180_ (.A1(\output_c[6][28] ),
    .A2(_1618_),
    .B1(net387),
    .Y(_1620_));
 sky130_fd_sc_hd__nor2_1 _3181_ (.A(_1619_),
    .B(net388),
    .Y(_0807_));
 sky130_fd_sc_hd__xor2_1 _3182_ (.A(net412),
    .B(_1618_),
    .X(_0806_));
 sky130_fd_sc_hd__buf_1 _3183_ (.A(\output_c[6][24] ),
    .X(_1621_));
 sky130_fd_sc_hd__and3_1 _3184_ (.A(_1604_),
    .B(_1607_),
    .C(_1617_),
    .X(_1622_));
 sky130_fd_sc_hd__a41o_1 _3185_ (.A1(\output_c[6][26] ),
    .A2(\output_c[6][25] ),
    .A3(_1621_),
    .A4(_1622_),
    .B1(\output_c[6][27] ),
    .X(_1623_));
 sky130_fd_sc_hd__and2b_1 _3186_ (.A_N(_1618_),
    .B(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__clkbuf_1 _3187_ (.A(_1624_),
    .X(_0805_));
 sky130_fd_sc_hd__buf_1 _3188_ (.A(_1622_),
    .X(_1625_));
 sky130_fd_sc_hd__nand3_1 _3189_ (.A(\output_c[6][25] ),
    .B(_1621_),
    .C(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__xnor2_1 _3190_ (.A(net213),
    .B(_1626_),
    .Y(_0804_));
 sky130_fd_sc_hd__a21o_1 _3191_ (.A1(_1621_),
    .A2(_1625_),
    .B1(\output_c[6][25] ),
    .X(_1627_));
 sky130_fd_sc_hd__and2_1 _3192_ (.A(_1626_),
    .B(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__clkbuf_1 _3193_ (.A(_1628_),
    .X(_0803_));
 sky130_fd_sc_hd__xor2_1 _3194_ (.A(_1621_),
    .B(_1625_),
    .X(_0802_));
 sky130_fd_sc_hd__buf_1 _3195_ (.A(_1607_),
    .X(_1629_));
 sky130_fd_sc_hd__a41o_1 _3196_ (.A1(\output_c[6][22] ),
    .A2(_1603_),
    .A3(_1629_),
    .A4(_1613_),
    .B1(\output_c[6][23] ),
    .X(_1630_));
 sky130_fd_sc_hd__and2b_1 _3197_ (.A_N(_1625_),
    .B(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _3198_ (.A(_1631_),
    .X(_0801_));
 sky130_fd_sc_hd__buf_1 _3199_ (.A(_1617_),
    .X(_1632_));
 sky130_fd_sc_hd__and3_1 _3200_ (.A(_1602_),
    .B(_1629_),
    .C(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__and3_1 _3201_ (.A(\output_c[6][21] ),
    .B(\output_c[6][20] ),
    .C(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__xor2_1 _3202_ (.A(net125),
    .B(_1634_),
    .X(_0800_));
 sky130_fd_sc_hd__a21oi_1 _3203_ (.A1(\output_c[6][20] ),
    .A2(_1633_),
    .B1(net243),
    .Y(_1635_));
 sky130_fd_sc_hd__nor2_1 _3204_ (.A(_1634_),
    .B(net244),
    .Y(_0799_));
 sky130_fd_sc_hd__xor2_1 _3205_ (.A(net299),
    .B(_1633_),
    .X(_0798_));
 sky130_fd_sc_hd__and3_1 _3206_ (.A(\output_c[6][16] ),
    .B(_1629_),
    .C(_1632_),
    .X(_1636_));
 sky130_fd_sc_hd__and3_1 _3207_ (.A(\output_c[6][18] ),
    .B(\output_c[6][17] ),
    .C(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__o21ba_1 _3208_ (.A1(net123),
    .A2(_1637_),
    .B1_N(_1633_),
    .X(_0797_));
 sky130_fd_sc_hd__a21oi_1 _3209_ (.A1(\output_c[6][17] ),
    .A2(_1636_),
    .B1(net228),
    .Y(_1638_));
 sky130_fd_sc_hd__nor2_1 _3210_ (.A(_1637_),
    .B(net229),
    .Y(_0796_));
 sky130_fd_sc_hd__xor2_1 _3211_ (.A(net301),
    .B(_1636_),
    .X(_0795_));
 sky130_fd_sc_hd__buf_1 _3212_ (.A(_1632_),
    .X(_1639_));
 sky130_fd_sc_hd__a21o_1 _3213_ (.A1(_1629_),
    .A2(_1639_),
    .B1(\output_c[6][16] ),
    .X(_1640_));
 sky130_fd_sc_hd__and2b_1 _3214_ (.A_N(_1636_),
    .B(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__clkbuf_1 _3215_ (.A(_1641_),
    .X(_0794_));
 sky130_fd_sc_hd__and3_1 _3216_ (.A(\output_c[6][12] ),
    .B(_1605_),
    .C(_1613_),
    .X(_1642_));
 sky130_fd_sc_hd__and3_1 _3217_ (.A(\output_c[6][14] ),
    .B(\output_c[6][13] ),
    .C(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__xor2_1 _3218_ (.A(net55),
    .B(_1643_),
    .X(_0793_));
 sky130_fd_sc_hd__buf_1 _3219_ (.A(_1639_),
    .X(_1644_));
 sky130_fd_sc_hd__a21oi_1 _3220_ (.A1(_1606_),
    .A2(_1644_),
    .B1(net398),
    .Y(_1645_));
 sky130_fd_sc_hd__nor2_1 _3221_ (.A(_1643_),
    .B(_1645_),
    .Y(_0792_));
 sky130_fd_sc_hd__nor2_1 _3222_ (.A(net323),
    .B(_1642_),
    .Y(_1646_));
 sky130_fd_sc_hd__a21oi_1 _3223_ (.A1(_1606_),
    .A2(_1644_),
    .B1(_1646_),
    .Y(_0791_));
 sky130_fd_sc_hd__and2_1 _3224_ (.A(_1605_),
    .B(_1639_),
    .X(_1647_));
 sky130_fd_sc_hd__nor2_1 _3225_ (.A(net392),
    .B(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__nor2_1 _3226_ (.A(_1642_),
    .B(_1648_),
    .Y(_0790_));
 sky130_fd_sc_hd__and3_1 _3227_ (.A(\output_c[6][9] ),
    .B(\output_c[6][8] ),
    .C(_1632_),
    .X(_1649_));
 sky130_fd_sc_hd__a21oi_1 _3228_ (.A1(\output_c[6][10] ),
    .A2(_1649_),
    .B1(net102),
    .Y(_1650_));
 sky130_fd_sc_hd__nor2_1 _3229_ (.A(_1647_),
    .B(net103),
    .Y(_0789_));
 sky130_fd_sc_hd__xor2_1 _3230_ (.A(net139),
    .B(_1649_),
    .X(_0788_));
 sky130_fd_sc_hd__a21oi_1 _3231_ (.A1(net239),
    .A2(_1644_),
    .B1(net355),
    .Y(_1651_));
 sky130_fd_sc_hd__nor2_1 _3232_ (.A(_1649_),
    .B(_1651_),
    .Y(_0787_));
 sky130_fd_sc_hd__xor2_1 _3233_ (.A(net239),
    .B(_1644_),
    .X(_0786_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3234_ (.A(_1611_),
    .X(_1652_));
 sky130_fd_sc_hd__and3_1 _3235_ (.A(\output_c[6][5] ),
    .B(_1608_),
    .C(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__a21o_1 _3236_ (.A1(\output_c[6][6] ),
    .A2(_1653_),
    .B1(\output_c[6][7] ),
    .X(_1654_));
 sky130_fd_sc_hd__and2b_1 _3237_ (.A_N(_1639_),
    .B(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _3238_ (.A(_1655_),
    .X(_0785_));
 sky130_fd_sc_hd__xor2_1 _3239_ (.A(net274),
    .B(_1653_),
    .X(_0784_));
 sky130_fd_sc_hd__a21oi_1 _3240_ (.A1(_1608_),
    .A2(_1652_),
    .B1(net456),
    .Y(_1656_));
 sky130_fd_sc_hd__nor2_1 _3241_ (.A(_1653_),
    .B(_1656_),
    .Y(_0783_));
 sky130_fd_sc_hd__xor2_1 _3242_ (.A(_1608_),
    .B(_1652_),
    .X(_0782_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3243_ (.A(_1154_),
    .X(_1657_));
 sky130_fd_sc_hd__and3_1 _3244_ (.A(\output_c[6][1] ),
    .B(_1657_),
    .C(_1609_),
    .X(_1658_));
 sky130_fd_sc_hd__and2_1 _3245_ (.A(\output_c[6][2] ),
    .B(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__o21ba_1 _3246_ (.A1(net286),
    .A2(_1659_),
    .B1_N(_1652_),
    .X(_0781_));
 sky130_fd_sc_hd__nor2_1 _3247_ (.A(net450),
    .B(_1658_),
    .Y(_1660_));
 sky130_fd_sc_hd__nor2_1 _3248_ (.A(_1659_),
    .B(_1660_),
    .Y(_0780_));
 sky130_fd_sc_hd__a21oi_1 _3249_ (.A1(_1597_),
    .A2(_1609_),
    .B1(net367),
    .Y(_1661_));
 sky130_fd_sc_hd__nor2_1 _3250_ (.A(_1658_),
    .B(_1661_),
    .Y(_0779_));
 sky130_fd_sc_hd__buf_1 _3251_ (.A(_1147_),
    .X(_1662_));
 sky130_fd_sc_hd__buf_1 _3252_ (.A(_1155_),
    .X(_1663_));
 sky130_fd_sc_hd__and3_1 _3253_ (.A(_1599_),
    .B(\input_a[6][0] ),
    .C(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__o2bb2a_1 _3254_ (.A1_N(_1662_),
    .A2_N(_1609_),
    .B1(_1664_),
    .B2(net191),
    .X(_0778_));
 sky130_fd_sc_hd__and4_1 _3255_ (.A(\output_c[5][27] ),
    .B(\output_c[5][26] ),
    .C(\output_c[5][25] ),
    .D(\output_c[5][24] ),
    .X(_1665_));
 sky130_fd_sc_hd__and4_1 _3256_ (.A(\output_c[5][19] ),
    .B(\output_c[5][18] ),
    .C(\output_c[5][17] ),
    .D(\output_c[5][16] ),
    .X(_1666_));
 sky130_fd_sc_hd__and3_1 _3257_ (.A(\output_c[5][21] ),
    .B(\output_c[5][20] ),
    .C(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__and3_1 _3258_ (.A(\output_c[5][23] ),
    .B(\output_c[5][22] ),
    .C(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__and4_1 _3259_ (.A(\output_c[5][11] ),
    .B(\output_c[5][10] ),
    .C(\output_c[5][9] ),
    .D(\output_c[5][8] ),
    .X(_1669_));
 sky130_fd_sc_hd__and3_1 _3260_ (.A(\output_c[5][13] ),
    .B(\output_c[5][12] ),
    .C(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__and3_1 _3261_ (.A(\output_c[5][15] ),
    .B(\output_c[5][14] ),
    .C(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__buf_1 _3262_ (.A(\output_c[5][4] ),
    .X(_1672_));
 sky130_fd_sc_hd__and3_1 _3263_ (.A(\output_c[5][0] ),
    .B(_1424_),
    .C(\input_a[5][0] ),
    .X(_1673_));
 sky130_fd_sc_hd__and2_1 _3264_ (.A(\output_c[5][3] ),
    .B(\output_c[5][2] ),
    .X(_1674_));
 sky130_fd_sc_hd__and4_1 _3265_ (.A(\output_c[5][1] ),
    .B(_1288_),
    .C(_1673_),
    .D(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__and2_1 _3266_ (.A(\output_c[5][7] ),
    .B(\output_c[5][6] ),
    .X(_1676_));
 sky130_fd_sc_hd__and4_1 _3267_ (.A(\output_c[5][5] ),
    .B(_1672_),
    .C(_1675_),
    .D(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__and4_1 _3268_ (.A(_1665_),
    .B(_1668_),
    .C(_1671_),
    .D(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__and4_1 _3269_ (.A(\output_c[5][30] ),
    .B(\output_c[5][29] ),
    .C(net491),
    .D(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__xor2_1 _3270_ (.A(net47),
    .B(_1679_),
    .X(_0777_));
 sky130_fd_sc_hd__and2_1 _3271_ (.A(\output_c[5][6] ),
    .B(\output_c[5][5] ),
    .X(_1680_));
 sky130_fd_sc_hd__and4_1 _3272_ (.A(\output_c[5][7] ),
    .B(\output_c[5][4] ),
    .C(_1675_),
    .D(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__and4_1 _3273_ (.A(_1665_),
    .B(_1668_),
    .C(_1671_),
    .D(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__and3_1 _3274_ (.A(\output_c[5][29] ),
    .B(net491),
    .C(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__xor2_1 _3275_ (.A(net84),
    .B(_1683_),
    .X(_0776_));
 sky130_fd_sc_hd__a21oi_1 _3276_ (.A1(net312),
    .A2(_1682_),
    .B1(net316),
    .Y(_1684_));
 sky130_fd_sc_hd__nor2_1 _3277_ (.A(_1683_),
    .B(_1684_),
    .Y(_0775_));
 sky130_fd_sc_hd__xor2_1 _3278_ (.A(net312),
    .B(_1682_),
    .X(_0774_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3279_ (.A(\output_c[5][24] ),
    .X(_1685_));
 sky130_fd_sc_hd__and3_1 _3280_ (.A(_1668_),
    .B(_1671_),
    .C(_1681_),
    .X(_1686_));
 sky130_fd_sc_hd__a41o_1 _3281_ (.A1(\output_c[5][26] ),
    .A2(\output_c[5][25] ),
    .A3(_1685_),
    .A4(_1686_),
    .B1(\output_c[5][27] ),
    .X(_1687_));
 sky130_fd_sc_hd__and2b_1 _3282_ (.A_N(_1682_),
    .B(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__clkbuf_1 _3283_ (.A(_1688_),
    .X(_0773_));
 sky130_fd_sc_hd__buf_1 _3284_ (.A(_1686_),
    .X(_1689_));
 sky130_fd_sc_hd__nand3_1 _3285_ (.A(\output_c[5][25] ),
    .B(_1685_),
    .C(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__xnor2_1 _3286_ (.A(net231),
    .B(_1690_),
    .Y(_0772_));
 sky130_fd_sc_hd__a21o_1 _3287_ (.A1(_1685_),
    .A2(_1689_),
    .B1(\output_c[5][25] ),
    .X(_1691_));
 sky130_fd_sc_hd__and2_1 _3288_ (.A(_1690_),
    .B(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__clkbuf_1 _3289_ (.A(_1692_),
    .X(_0771_));
 sky130_fd_sc_hd__xor2_1 _3290_ (.A(_1685_),
    .B(_1689_),
    .X(_0770_));
 sky130_fd_sc_hd__buf_1 _3291_ (.A(_1671_),
    .X(_1693_));
 sky130_fd_sc_hd__a41o_1 _3292_ (.A1(\output_c[5][22] ),
    .A2(_1667_),
    .A3(_1693_),
    .A4(_1677_),
    .B1(\output_c[5][23] ),
    .X(_1694_));
 sky130_fd_sc_hd__and2b_1 _3293_ (.A_N(_1689_),
    .B(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _3294_ (.A(_1695_),
    .X(_0769_));
 sky130_fd_sc_hd__buf_1 _3295_ (.A(_1681_),
    .X(_1696_));
 sky130_fd_sc_hd__and3_1 _3296_ (.A(_1666_),
    .B(_1693_),
    .C(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__and3_1 _3297_ (.A(\output_c[5][21] ),
    .B(\output_c[5][20] ),
    .C(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__xor2_1 _3298_ (.A(net152),
    .B(_1698_),
    .X(_0768_));
 sky130_fd_sc_hd__a21oi_1 _3299_ (.A1(net314),
    .A2(_1697_),
    .B1(net417),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_1 _3300_ (.A(_1698_),
    .B(_1699_),
    .Y(_0767_));
 sky130_fd_sc_hd__xor2_1 _3301_ (.A(net314),
    .B(_1697_),
    .X(_0766_));
 sky130_fd_sc_hd__and3_1 _3302_ (.A(\output_c[5][16] ),
    .B(_1693_),
    .C(_1696_),
    .X(_1700_));
 sky130_fd_sc_hd__and3_1 _3303_ (.A(\output_c[5][18] ),
    .B(\output_c[5][17] ),
    .C(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__o21ba_1 _3304_ (.A1(net223),
    .A2(_1701_),
    .B1_N(_1697_),
    .X(_0765_));
 sky130_fd_sc_hd__a21oi_1 _3305_ (.A1(net386),
    .A2(_1700_),
    .B1(net423),
    .Y(_1702_));
 sky130_fd_sc_hd__nor2_1 _3306_ (.A(_1701_),
    .B(_1702_),
    .Y(_0764_));
 sky130_fd_sc_hd__xor2_1 _3307_ (.A(net386),
    .B(_1700_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_1 _3308_ (.A(_1696_),
    .X(_1703_));
 sky130_fd_sc_hd__a21o_1 _3309_ (.A1(_1693_),
    .A2(_1703_),
    .B1(\output_c[5][16] ),
    .X(_1704_));
 sky130_fd_sc_hd__and2b_1 _3310_ (.A_N(_1700_),
    .B(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__clkbuf_1 _3311_ (.A(_1705_),
    .X(_0762_));
 sky130_fd_sc_hd__and3_1 _3312_ (.A(\output_c[5][12] ),
    .B(_1669_),
    .C(_1677_),
    .X(_1706_));
 sky130_fd_sc_hd__and3_1 _3313_ (.A(\output_c[5][14] ),
    .B(\output_c[5][13] ),
    .C(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__xor2_1 _3314_ (.A(net61),
    .B(_1707_),
    .X(_0761_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3315_ (.A(_1703_),
    .X(_1708_));
 sky130_fd_sc_hd__a21oi_1 _3316_ (.A1(_1670_),
    .A2(_1708_),
    .B1(net224),
    .Y(_1709_));
 sky130_fd_sc_hd__nor2_1 _3317_ (.A(_1707_),
    .B(_1709_),
    .Y(_0760_));
 sky130_fd_sc_hd__nor2_1 _3318_ (.A(net340),
    .B(_1706_),
    .Y(_1710_));
 sky130_fd_sc_hd__a21oi_1 _3319_ (.A1(_1670_),
    .A2(_1708_),
    .B1(_1710_),
    .Y(_0759_));
 sky130_fd_sc_hd__and2_1 _3320_ (.A(_1669_),
    .B(_1703_),
    .X(_1711_));
 sky130_fd_sc_hd__nor2_1 _3321_ (.A(net459),
    .B(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__nor2_1 _3322_ (.A(_1706_),
    .B(_1712_),
    .Y(_0758_));
 sky130_fd_sc_hd__and3_1 _3323_ (.A(\output_c[5][9] ),
    .B(\output_c[5][8] ),
    .C(_1696_),
    .X(_1713_));
 sky130_fd_sc_hd__a21oi_1 _3324_ (.A1(net121),
    .A2(_1713_),
    .B1(net133),
    .Y(_1714_));
 sky130_fd_sc_hd__nor2_1 _3325_ (.A(_1711_),
    .B(_1714_),
    .Y(_0757_));
 sky130_fd_sc_hd__xor2_1 _3326_ (.A(net121),
    .B(_1713_),
    .X(_0756_));
 sky130_fd_sc_hd__a21oi_1 _3327_ (.A1(\output_c[5][8] ),
    .A2(_1708_),
    .B1(net187),
    .Y(_1715_));
 sky130_fd_sc_hd__nor2_1 _3328_ (.A(_1713_),
    .B(net188),
    .Y(_0755_));
 sky130_fd_sc_hd__xor2_1 _3329_ (.A(net250),
    .B(_1708_),
    .X(_0754_));
 sky130_fd_sc_hd__buf_1 _3330_ (.A(_1675_),
    .X(_1716_));
 sky130_fd_sc_hd__and3_1 _3331_ (.A(\output_c[5][5] ),
    .B(_1672_),
    .C(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__a21o_1 _3332_ (.A1(\output_c[5][6] ),
    .A2(_1717_),
    .B1(\output_c[5][7] ),
    .X(_1718_));
 sky130_fd_sc_hd__and2b_1 _3333_ (.A_N(_1703_),
    .B(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_1 _3334_ (.A(_1719_),
    .X(_0753_));
 sky130_fd_sc_hd__xor2_1 _3335_ (.A(net365),
    .B(_1717_),
    .X(_0752_));
 sky130_fd_sc_hd__a21oi_1 _3336_ (.A1(_1672_),
    .A2(_1716_),
    .B1(net471),
    .Y(_1720_));
 sky130_fd_sc_hd__nor2_1 _3337_ (.A(_1717_),
    .B(_1720_),
    .Y(_0751_));
 sky130_fd_sc_hd__xor2_1 _3338_ (.A(_1672_),
    .B(_1716_),
    .X(_0750_));
 sky130_fd_sc_hd__and3_1 _3339_ (.A(\output_c[5][1] ),
    .B(_1657_),
    .C(_1673_),
    .X(_1721_));
 sky130_fd_sc_hd__and2_1 _3340_ (.A(\output_c[5][2] ),
    .B(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__o21ba_1 _3341_ (.A1(net371),
    .A2(_1722_),
    .B1_N(_1716_),
    .X(_0749_));
 sky130_fd_sc_hd__nor2_1 _3342_ (.A(net440),
    .B(_1721_),
    .Y(_1723_));
 sky130_fd_sc_hd__nor2_1 _3343_ (.A(_1722_),
    .B(_1723_),
    .Y(_0748_));
 sky130_fd_sc_hd__a21oi_1 _3344_ (.A1(_1597_),
    .A2(_1673_),
    .B1(net348),
    .Y(_1724_));
 sky130_fd_sc_hd__nor2_1 _3345_ (.A(_1721_),
    .B(_1724_),
    .Y(_0747_));
 sky130_fd_sc_hd__and3_1 _3346_ (.A(_1599_),
    .B(\input_a[5][0] ),
    .C(_1663_),
    .X(_1725_));
 sky130_fd_sc_hd__o2bb2a_1 _3347_ (.A1_N(_1662_),
    .A2_N(_1673_),
    .B1(_1725_),
    .B2(net180),
    .X(_0746_));
 sky130_fd_sc_hd__and4_1 _3348_ (.A(\output_c[4][27] ),
    .B(\output_c[4][26] ),
    .C(\output_c[4][25] ),
    .D(\output_c[4][24] ),
    .X(_1726_));
 sky130_fd_sc_hd__and4_1 _3349_ (.A(\output_c[4][11] ),
    .B(\output_c[4][10] ),
    .C(\output_c[4][9] ),
    .D(\output_c[4][8] ),
    .X(_1727_));
 sky130_fd_sc_hd__and3_1 _3350_ (.A(\output_c[4][13] ),
    .B(\output_c[4][12] ),
    .C(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__and3_1 _3351_ (.A(\output_c[4][15] ),
    .B(\output_c[4][14] ),
    .C(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__buf_1 _3352_ (.A(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__buf_1 _3353_ (.A(\output_c[4][4] ),
    .X(_1731_));
 sky130_fd_sc_hd__and3_1 _3354_ (.A(\output_c[4][0] ),
    .B(_1070_),
    .C(\input_a[4][0] ),
    .X(_1732_));
 sky130_fd_sc_hd__and2_1 _3355_ (.A(\output_c[4][3] ),
    .B(\output_c[4][2] ),
    .X(_1733_));
 sky130_fd_sc_hd__and4_1 _3356_ (.A(\output_c[4][1] ),
    .B(_1164_),
    .C(_1732_),
    .D(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__and2_1 _3357_ (.A(\output_c[4][7] ),
    .B(\output_c[4][6] ),
    .X(_1735_));
 sky130_fd_sc_hd__and4_1 _3358_ (.A(\output_c[4][5] ),
    .B(_1731_),
    .C(_1734_),
    .D(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__and2_1 _3359_ (.A(\output_c[4][21] ),
    .B(\output_c[4][20] ),
    .X(_1737_));
 sky130_fd_sc_hd__and4_1 _3360_ (.A(\output_c[4][19] ),
    .B(\output_c[4][18] ),
    .C(\output_c[4][17] ),
    .D(\output_c[4][16] ),
    .X(_1738_));
 sky130_fd_sc_hd__and4_1 _3361_ (.A(\output_c[4][23] ),
    .B(\output_c[4][22] ),
    .C(_1737_),
    .D(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__and4_1 _3362_ (.A(_1726_),
    .B(_1730_),
    .C(_1736_),
    .D(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__and4_1 _3363_ (.A(\output_c[4][30] ),
    .B(\output_c[4][29] ),
    .C(\output_c[4][28] ),
    .D(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__xor2_1 _3364_ (.A(net38),
    .B(_1741_),
    .X(_0745_));
 sky130_fd_sc_hd__and2_1 _3365_ (.A(\output_c[4][6] ),
    .B(\output_c[4][5] ),
    .X(_1742_));
 sky130_fd_sc_hd__and4_1 _3366_ (.A(\output_c[4][7] ),
    .B(\output_c[4][4] ),
    .C(_1734_),
    .D(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__and4_1 _3367_ (.A(\output_c[4][23] ),
    .B(\output_c[4][22] ),
    .C(_1737_),
    .D(_1738_),
    .X(_1744_));
 sky130_fd_sc_hd__and3_1 _3368_ (.A(_1729_),
    .B(_1743_),
    .C(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__and4_1 _3369_ (.A(\output_c[4][29] ),
    .B(\output_c[4][28] ),
    .C(_1726_),
    .D(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__xor2_1 _3370_ (.A(net81),
    .B(_1746_),
    .X(_0744_));
 sky130_fd_sc_hd__a21oi_1 _3371_ (.A1(\output_c[4][28] ),
    .A2(_1740_),
    .B1(net362),
    .Y(_1747_));
 sky130_fd_sc_hd__nor2_1 _3372_ (.A(_1746_),
    .B(net363),
    .Y(_0743_));
 sky130_fd_sc_hd__xor2_1 _3373_ (.A(net368),
    .B(_1740_),
    .X(_0742_));
 sky130_fd_sc_hd__buf_1 _3374_ (.A(\output_c[4][24] ),
    .X(_1748_));
 sky130_fd_sc_hd__a41o_1 _3375_ (.A1(\output_c[4][26] ),
    .A2(\output_c[4][25] ),
    .A3(_1748_),
    .A4(_1745_),
    .B1(\output_c[4][27] ),
    .X(_1749_));
 sky130_fd_sc_hd__and2b_1 _3376_ (.A_N(_1740_),
    .B(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__clkbuf_1 _3377_ (.A(_1750_),
    .X(_0741_));
 sky130_fd_sc_hd__buf_1 _3378_ (.A(_1745_),
    .X(_1751_));
 sky130_fd_sc_hd__and3_1 _3379_ (.A(\output_c[4][25] ),
    .B(_1748_),
    .C(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__xor2_1 _3380_ (.A(net120),
    .B(_1752_),
    .X(_0740_));
 sky130_fd_sc_hd__a21oi_1 _3381_ (.A1(_1748_),
    .A2(_1751_),
    .B1(net474),
    .Y(_1753_));
 sky130_fd_sc_hd__nor2_1 _3382_ (.A(_1752_),
    .B(_1753_),
    .Y(_0739_));
 sky130_fd_sc_hd__xor2_1 _3383_ (.A(_1748_),
    .B(_1751_),
    .X(_0738_));
 sky130_fd_sc_hd__buf_1 _3384_ (.A(_1743_),
    .X(_1754_));
 sky130_fd_sc_hd__and3_1 _3385_ (.A(_1729_),
    .B(_1738_),
    .C(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__buf_1 _3386_ (.A(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__and3_1 _3387_ (.A(\output_c[4][22] ),
    .B(_1737_),
    .C(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__o21ba_1 _3388_ (.A1(net402),
    .A2(_1757_),
    .B1_N(_1751_),
    .X(_0737_));
 sky130_fd_sc_hd__and2_1 _3389_ (.A(_1737_),
    .B(_1755_),
    .X(_1758_));
 sky130_fd_sc_hd__xor2_1 _3390_ (.A(net366),
    .B(_1758_),
    .X(_0736_));
 sky130_fd_sc_hd__a21oi_1 _3391_ (.A1(net114),
    .A2(_1756_),
    .B1(net131),
    .Y(_1759_));
 sky130_fd_sc_hd__nor2_1 _3392_ (.A(_1758_),
    .B(_1759_),
    .Y(_0735_));
 sky130_fd_sc_hd__xor2_1 _3393_ (.A(net114),
    .B(_1756_),
    .X(_0734_));
 sky130_fd_sc_hd__and4_1 _3394_ (.A(\output_c[4][17] ),
    .B(\output_c[4][16] ),
    .C(_1730_),
    .D(_1736_),
    .X(_1760_));
 sky130_fd_sc_hd__a21o_1 _3395_ (.A1(\output_c[4][18] ),
    .A2(_1760_),
    .B1(\output_c[4][19] ),
    .X(_1761_));
 sky130_fd_sc_hd__and2b_1 _3396_ (.A_N(_1756_),
    .B(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__clkbuf_1 _3397_ (.A(_1762_),
    .X(_0733_));
 sky130_fd_sc_hd__xor2_1 _3398_ (.A(net190),
    .B(_1760_),
    .X(_0732_));
 sky130_fd_sc_hd__and3_1 _3399_ (.A(\output_c[4][16] ),
    .B(_1730_),
    .C(_1754_),
    .X(_1763_));
 sky130_fd_sc_hd__nor2_1 _3400_ (.A(net397),
    .B(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__nor2_1 _3401_ (.A(_1760_),
    .B(_1764_),
    .Y(_0731_));
 sky130_fd_sc_hd__buf_1 _3402_ (.A(_1754_),
    .X(_1765_));
 sky130_fd_sc_hd__buf_1 _3403_ (.A(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__a21oi_1 _3404_ (.A1(_1730_),
    .A2(_1766_),
    .B1(net444),
    .Y(_1767_));
 sky130_fd_sc_hd__nor2_1 _3405_ (.A(_1763_),
    .B(_1767_),
    .Y(_0730_));
 sky130_fd_sc_hd__and3_1 _3406_ (.A(\output_c[4][12] ),
    .B(_1727_),
    .C(_1736_),
    .X(_1768_));
 sky130_fd_sc_hd__and3_1 _3407_ (.A(\output_c[4][14] ),
    .B(\output_c[4][13] ),
    .C(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__xor2_1 _3408_ (.A(net65),
    .B(_1769_),
    .X(_0729_));
 sky130_fd_sc_hd__a21oi_1 _3409_ (.A1(_1728_),
    .A2(_1766_),
    .B1(net373),
    .Y(_1770_));
 sky130_fd_sc_hd__nor2_1 _3410_ (.A(_1769_),
    .B(_1770_),
    .Y(_0728_));
 sky130_fd_sc_hd__nor2_1 _3411_ (.A(net240),
    .B(_1768_),
    .Y(_1771_));
 sky130_fd_sc_hd__a21oi_1 _3412_ (.A1(_1728_),
    .A2(_1766_),
    .B1(_1771_),
    .Y(_0727_));
 sky130_fd_sc_hd__and2_1 _3413_ (.A(_1727_),
    .B(_1765_),
    .X(_1772_));
 sky130_fd_sc_hd__nor2_1 _3414_ (.A(net457),
    .B(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__nor2_1 _3415_ (.A(_1768_),
    .B(_1773_),
    .Y(_0726_));
 sky130_fd_sc_hd__and3_1 _3416_ (.A(\output_c[4][9] ),
    .B(\output_c[4][8] ),
    .C(_1754_),
    .X(_1774_));
 sky130_fd_sc_hd__a21oi_1 _3417_ (.A1(net106),
    .A2(_1774_),
    .B1(net111),
    .Y(_1775_));
 sky130_fd_sc_hd__nor2_1 _3418_ (.A(_1772_),
    .B(_1775_),
    .Y(_0725_));
 sky130_fd_sc_hd__xor2_1 _3419_ (.A(net106),
    .B(_1774_),
    .X(_0724_));
 sky130_fd_sc_hd__a21oi_1 _3420_ (.A1(\output_c[4][8] ),
    .A2(_1765_),
    .B1(net302),
    .Y(_1776_));
 sky130_fd_sc_hd__nor2_1 _3421_ (.A(_1774_),
    .B(net303),
    .Y(_0723_));
 sky130_fd_sc_hd__xor2_1 _3422_ (.A(net315),
    .B(_1766_),
    .X(_0722_));
 sky130_fd_sc_hd__buf_1 _3423_ (.A(_1734_),
    .X(_1777_));
 sky130_fd_sc_hd__and3_1 _3424_ (.A(\output_c[4][5] ),
    .B(_1731_),
    .C(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__a21o_1 _3425_ (.A1(\output_c[4][6] ),
    .A2(_1778_),
    .B1(\output_c[4][7] ),
    .X(_1779_));
 sky130_fd_sc_hd__and2b_1 _3426_ (.A_N(_1765_),
    .B(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__clkbuf_1 _3427_ (.A(_1780_),
    .X(_0721_));
 sky130_fd_sc_hd__xor2_1 _3428_ (.A(net324),
    .B(_1778_),
    .X(_0720_));
 sky130_fd_sc_hd__a21oi_1 _3429_ (.A1(_1731_),
    .A2(_1777_),
    .B1(net468),
    .Y(_1781_));
 sky130_fd_sc_hd__nor2_1 _3430_ (.A(_1778_),
    .B(_1781_),
    .Y(_0719_));
 sky130_fd_sc_hd__xor2_1 _3431_ (.A(_1731_),
    .B(_1777_),
    .X(_0718_));
 sky130_fd_sc_hd__and3_1 _3432_ (.A(\output_c[4][1] ),
    .B(_1657_),
    .C(_1732_),
    .X(_1782_));
 sky130_fd_sc_hd__and2_1 _3433_ (.A(\output_c[4][2] ),
    .B(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__o21ba_1 _3434_ (.A1(net289),
    .A2(_1783_),
    .B1_N(_1777_),
    .X(_0717_));
 sky130_fd_sc_hd__nor2_1 _3435_ (.A(net438),
    .B(_1782_),
    .Y(_1784_));
 sky130_fd_sc_hd__nor2_1 _3436_ (.A(_1783_),
    .B(_1784_),
    .Y(_0716_));
 sky130_fd_sc_hd__a21oi_1 _3437_ (.A1(_1597_),
    .A2(_1732_),
    .B1(net207),
    .Y(_1785_));
 sky130_fd_sc_hd__nor2_1 _3438_ (.A(_1782_),
    .B(_1785_),
    .Y(_0715_));
 sky130_fd_sc_hd__and3_1 _3439_ (.A(_1599_),
    .B(\input_a[4][0] ),
    .C(_1663_),
    .X(_1786_));
 sky130_fd_sc_hd__o2bb2a_1 _3440_ (.A1_N(_1662_),
    .A2_N(_1732_),
    .B1(_1786_),
    .B2(net233),
    .X(_0714_));
 sky130_fd_sc_hd__and4_1 _3441_ (.A(\output_c[3][27] ),
    .B(\output_c[3][26] ),
    .C(\output_c[3][25] ),
    .D(\output_c[3][24] ),
    .X(_1787_));
 sky130_fd_sc_hd__and4_1 _3442_ (.A(\output_c[3][19] ),
    .B(\output_c[3][18] ),
    .C(\output_c[3][17] ),
    .D(\output_c[3][16] ),
    .X(_1788_));
 sky130_fd_sc_hd__and3_1 _3443_ (.A(\output_c[3][21] ),
    .B(\output_c[3][20] ),
    .C(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__and3_1 _3444_ (.A(\output_c[3][23] ),
    .B(\output_c[3][22] ),
    .C(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__and4_1 _3445_ (.A(\output_c[3][11] ),
    .B(\output_c[3][10] ),
    .C(\output_c[3][9] ),
    .D(\output_c[3][8] ),
    .X(_1791_));
 sky130_fd_sc_hd__and3_1 _3446_ (.A(\output_c[3][13] ),
    .B(\output_c[3][12] ),
    .C(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__and3_1 _3447_ (.A(\output_c[3][15] ),
    .B(\output_c[3][14] ),
    .C(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__and3_1 _3448_ (.A(\output_c[3][0] ),
    .B(_1289_),
    .C(\input_a[3][0] ),
    .X(_1794_));
 sky130_fd_sc_hd__and2_1 _3449_ (.A(\output_c[3][3] ),
    .B(\output_c[3][2] ),
    .X(_1795_));
 sky130_fd_sc_hd__and4_1 _3450_ (.A(\output_c[3][1] ),
    .B(_1288_),
    .C(_1794_),
    .D(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__and2_1 _3451_ (.A(\output_c[3][7] ),
    .B(\output_c[3][6] ),
    .X(_1797_));
 sky130_fd_sc_hd__and4_1 _3452_ (.A(\output_c[3][5] ),
    .B(\output_c[3][4] ),
    .C(_1796_),
    .D(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__and4_1 _3453_ (.A(_1787_),
    .B(_1790_),
    .C(_1793_),
    .D(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__and4_1 _3454_ (.A(\output_c[3][30] ),
    .B(\output_c[3][29] ),
    .C(\output_c[3][28] ),
    .D(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__xor2_1 _3455_ (.A(net45),
    .B(_1800_),
    .X(_0713_));
 sky130_fd_sc_hd__and2_1 _3456_ (.A(\output_c[3][6] ),
    .B(\output_c[3][5] ),
    .X(_1801_));
 sky130_fd_sc_hd__and4_1 _3457_ (.A(\output_c[3][7] ),
    .B(\output_c[3][4] ),
    .C(_1796_),
    .D(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__and4_1 _3458_ (.A(_1787_),
    .B(_1790_),
    .C(_1793_),
    .D(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__and3_1 _3459_ (.A(\output_c[3][29] ),
    .B(\output_c[3][28] ),
    .C(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__xor2_1 _3460_ (.A(net85),
    .B(_1804_),
    .X(_0712_));
 sky130_fd_sc_hd__a21oi_1 _3461_ (.A1(net256),
    .A2(_1803_),
    .B1(net263),
    .Y(_1805_));
 sky130_fd_sc_hd__nor2_1 _3462_ (.A(_1804_),
    .B(_1805_),
    .Y(_0711_));
 sky130_fd_sc_hd__xor2_1 _3463_ (.A(net256),
    .B(_1803_),
    .X(_0710_));
 sky130_fd_sc_hd__buf_1 _3464_ (.A(\output_c[3][24] ),
    .X(_1806_));
 sky130_fd_sc_hd__and3_1 _3465_ (.A(_1790_),
    .B(_1793_),
    .C(_1802_),
    .X(_1807_));
 sky130_fd_sc_hd__a41o_1 _3466_ (.A1(\output_c[3][26] ),
    .A2(\output_c[3][25] ),
    .A3(_1806_),
    .A4(_1807_),
    .B1(\output_c[3][27] ),
    .X(_1808_));
 sky130_fd_sc_hd__and2b_1 _3467_ (.A_N(_1803_),
    .B(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__clkbuf_1 _3468_ (.A(_1809_),
    .X(_0709_));
 sky130_fd_sc_hd__buf_1 _3469_ (.A(_1807_),
    .X(_1810_));
 sky130_fd_sc_hd__nand3_1 _3470_ (.A(\output_c[3][25] ),
    .B(_1806_),
    .C(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__xnor2_1 _3471_ (.A(net209),
    .B(_1811_),
    .Y(_0708_));
 sky130_fd_sc_hd__a21o_1 _3472_ (.A1(_1806_),
    .A2(_1810_),
    .B1(\output_c[3][25] ),
    .X(_1812_));
 sky130_fd_sc_hd__and2_1 _3473_ (.A(_1811_),
    .B(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _3474_ (.A(_1813_),
    .X(_0707_));
 sky130_fd_sc_hd__xor2_1 _3475_ (.A(_1806_),
    .B(_1810_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_1 _3476_ (.A(_1793_),
    .X(_1814_));
 sky130_fd_sc_hd__a41o_1 _3477_ (.A1(\output_c[3][22] ),
    .A2(_1789_),
    .A3(_1814_),
    .A4(_1798_),
    .B1(\output_c[3][23] ),
    .X(_1815_));
 sky130_fd_sc_hd__and2b_1 _3478_ (.A_N(_1810_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_1 _3479_ (.A(_1816_),
    .X(_0705_));
 sky130_fd_sc_hd__buf_1 _3480_ (.A(_1802_),
    .X(_1817_));
 sky130_fd_sc_hd__and3_1 _3481_ (.A(_1788_),
    .B(_1814_),
    .C(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__and3_1 _3482_ (.A(\output_c[3][21] ),
    .B(\output_c[3][20] ),
    .C(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__xor2_1 _3483_ (.A(net100),
    .B(_1819_),
    .X(_0704_));
 sky130_fd_sc_hd__a21oi_1 _3484_ (.A1(\output_c[3][20] ),
    .A2(_1818_),
    .B1(net195),
    .Y(_1820_));
 sky130_fd_sc_hd__nor2_1 _3485_ (.A(_1819_),
    .B(net196),
    .Y(_0703_));
 sky130_fd_sc_hd__xor2_1 _3486_ (.A(net258),
    .B(_1818_),
    .X(_0702_));
 sky130_fd_sc_hd__and3_1 _3487_ (.A(\output_c[3][16] ),
    .B(_1814_),
    .C(_1817_),
    .X(_1821_));
 sky130_fd_sc_hd__and3_1 _3488_ (.A(\output_c[3][18] ),
    .B(\output_c[3][17] ),
    .C(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__o21ba_1 _3489_ (.A1(net134),
    .A2(_1822_),
    .B1_N(_1818_),
    .X(_0701_));
 sky130_fd_sc_hd__a21oi_1 _3490_ (.A1(net278),
    .A2(_1821_),
    .B1(net322),
    .Y(_1823_));
 sky130_fd_sc_hd__nor2_1 _3491_ (.A(_1822_),
    .B(_1823_),
    .Y(_0700_));
 sky130_fd_sc_hd__xor2_1 _3492_ (.A(net278),
    .B(_1821_),
    .X(_0699_));
 sky130_fd_sc_hd__buf_1 _3493_ (.A(_1817_),
    .X(_1824_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3494_ (.A(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__a21oi_1 _3495_ (.A1(_1814_),
    .A2(_1825_),
    .B1(net242),
    .Y(_1826_));
 sky130_fd_sc_hd__nor2_1 _3496_ (.A(_1821_),
    .B(_1826_),
    .Y(_0698_));
 sky130_fd_sc_hd__and3_1 _3497_ (.A(\output_c[3][12] ),
    .B(_1791_),
    .C(_1798_),
    .X(_1827_));
 sky130_fd_sc_hd__and3_1 _3498_ (.A(\output_c[3][14] ),
    .B(\output_c[3][13] ),
    .C(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__xor2_1 _3499_ (.A(net52),
    .B(_1828_),
    .X(_0697_));
 sky130_fd_sc_hd__a21oi_1 _3500_ (.A1(_1792_),
    .A2(_1825_),
    .B1(net235),
    .Y(_1829_));
 sky130_fd_sc_hd__nor2_1 _3501_ (.A(_1828_),
    .B(_1829_),
    .Y(_0696_));
 sky130_fd_sc_hd__nor2_1 _3502_ (.A(net245),
    .B(_1827_),
    .Y(_1830_));
 sky130_fd_sc_hd__a21oi_1 _3503_ (.A1(_1792_),
    .A2(_1825_),
    .B1(_1830_),
    .Y(_0695_));
 sky130_fd_sc_hd__and2_1 _3504_ (.A(_1791_),
    .B(_1824_),
    .X(_1831_));
 sky130_fd_sc_hd__nor2_1 _3505_ (.A(net389),
    .B(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__nor2_1 _3506_ (.A(_1827_),
    .B(_1832_),
    .Y(_0694_));
 sky130_fd_sc_hd__and3_1 _3507_ (.A(\output_c[3][9] ),
    .B(\output_c[3][8] ),
    .C(_1817_),
    .X(_1833_));
 sky130_fd_sc_hd__a21oi_1 _3508_ (.A1(net92),
    .A2(_1833_),
    .B1(net179),
    .Y(_1834_));
 sky130_fd_sc_hd__nor2_1 _3509_ (.A(_1831_),
    .B(_1834_),
    .Y(_0693_));
 sky130_fd_sc_hd__xor2_1 _3510_ (.A(net92),
    .B(_1833_),
    .X(_0692_));
 sky130_fd_sc_hd__a21oi_1 _3511_ (.A1(net251),
    .A2(_1824_),
    .B1(net261),
    .Y(_1835_));
 sky130_fd_sc_hd__nor2_1 _3512_ (.A(_1833_),
    .B(_1835_),
    .Y(_0691_));
 sky130_fd_sc_hd__xor2_1 _3513_ (.A(net251),
    .B(_1825_),
    .X(_0690_));
 sky130_fd_sc_hd__buf_1 _3514_ (.A(\output_c[3][4] ),
    .X(_1836_));
 sky130_fd_sc_hd__a31o_1 _3515_ (.A1(_1836_),
    .A2(_1796_),
    .A3(_1801_),
    .B1(\output_c[3][7] ),
    .X(_1837_));
 sky130_fd_sc_hd__and2b_1 _3516_ (.A_N(_1824_),
    .B(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__clkbuf_1 _3517_ (.A(_1838_),
    .X(_0689_));
 sky130_fd_sc_hd__buf_1 _3518_ (.A(_1796_),
    .X(_1839_));
 sky130_fd_sc_hd__and3_1 _3519_ (.A(\output_c[3][5] ),
    .B(_1836_),
    .C(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__xor2_1 _3520_ (.A(net170),
    .B(_1840_),
    .X(_0688_));
 sky130_fd_sc_hd__a21oi_1 _3521_ (.A1(_1836_),
    .A2(_1839_),
    .B1(net482),
    .Y(_1841_));
 sky130_fd_sc_hd__nor2_1 _3522_ (.A(_1840_),
    .B(_1841_),
    .Y(_0687_));
 sky130_fd_sc_hd__xor2_1 _3523_ (.A(_1836_),
    .B(_1839_),
    .X(_0686_));
 sky130_fd_sc_hd__and3_1 _3524_ (.A(\output_c[3][1] ),
    .B(_1657_),
    .C(_1794_),
    .X(_1842_));
 sky130_fd_sc_hd__and2_1 _3525_ (.A(\output_c[3][2] ),
    .B(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__o21ba_1 _3526_ (.A1(net226),
    .A2(_1843_),
    .B1_N(_1839_),
    .X(_0685_));
 sky130_fd_sc_hd__nor2_1 _3527_ (.A(net445),
    .B(_1842_),
    .Y(_1844_));
 sky130_fd_sc_hd__nor2_1 _3528_ (.A(_1843_),
    .B(_1844_),
    .Y(_0684_));
 sky130_fd_sc_hd__clkbuf_2 _3529_ (.A(_1345_),
    .X(_1845_));
 sky130_fd_sc_hd__a21oi_1 _3530_ (.A1(_1845_),
    .A2(_1794_),
    .B1(net410),
    .Y(_1846_));
 sky130_fd_sc_hd__nor2_1 _3531_ (.A(_1842_),
    .B(_1846_),
    .Y(_0683_));
 sky130_fd_sc_hd__buf_1 _3532_ (.A(_1348_),
    .X(_1847_));
 sky130_fd_sc_hd__and3_1 _3533_ (.A(_1847_),
    .B(\input_a[3][0] ),
    .C(_1663_),
    .X(_1848_));
 sky130_fd_sc_hd__o2bb2a_1 _3534_ (.A1_N(_1662_),
    .A2_N(_1794_),
    .B1(_1848_),
    .B2(net183),
    .X(_0682_));
 sky130_fd_sc_hd__and4_1 _3535_ (.A(\output_c[2][27] ),
    .B(\output_c[2][26] ),
    .C(\output_c[2][25] ),
    .D(\output_c[2][24] ),
    .X(_1849_));
 sky130_fd_sc_hd__and4_1 _3536_ (.A(\output_c[2][19] ),
    .B(\output_c[2][18] ),
    .C(\output_c[2][17] ),
    .D(\output_c[2][16] ),
    .X(_1850_));
 sky130_fd_sc_hd__and3_1 _3537_ (.A(\output_c[2][21] ),
    .B(\output_c[2][20] ),
    .C(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__and3_1 _3538_ (.A(\output_c[2][23] ),
    .B(\output_c[2][22] ),
    .C(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__and4_1 _3539_ (.A(\output_c[2][11] ),
    .B(\output_c[2][10] ),
    .C(\output_c[2][9] ),
    .D(\output_c[2][8] ),
    .X(_1853_));
 sky130_fd_sc_hd__and3_1 _3540_ (.A(\output_c[2][13] ),
    .B(\output_c[2][12] ),
    .C(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__and3_1 _3541_ (.A(\output_c[2][15] ),
    .B(\output_c[2][14] ),
    .C(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__buf_1 _3542_ (.A(\output_c[2][4] ),
    .X(_1856_));
 sky130_fd_sc_hd__and3_1 _3543_ (.A(\output_c[2][0] ),
    .B(_1424_),
    .C(\input_a[2][0] ),
    .X(_1857_));
 sky130_fd_sc_hd__and2_1 _3544_ (.A(\output_c[2][3] ),
    .B(\output_c[2][2] ),
    .X(_1858_));
 sky130_fd_sc_hd__and4_1 _3545_ (.A(\output_c[2][1] ),
    .B(_1288_),
    .C(_1857_),
    .D(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__and2_1 _3546_ (.A(\output_c[2][7] ),
    .B(\output_c[2][6] ),
    .X(_1860_));
 sky130_fd_sc_hd__and4_1 _3547_ (.A(\output_c[2][5] ),
    .B(_1856_),
    .C(_1859_),
    .D(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__and4_1 _3548_ (.A(_1849_),
    .B(_1852_),
    .C(_1855_),
    .D(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__and4_1 _3549_ (.A(\output_c[2][30] ),
    .B(\output_c[2][29] ),
    .C(\output_c[2][28] ),
    .D(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__xor2_1 _3550_ (.A(net42),
    .B(_1863_),
    .X(_0681_));
 sky130_fd_sc_hd__and2_1 _3551_ (.A(\output_c[2][6] ),
    .B(\output_c[2][5] ),
    .X(_1864_));
 sky130_fd_sc_hd__and4_1 _3552_ (.A(\output_c[2][7] ),
    .B(\output_c[2][4] ),
    .C(_1859_),
    .D(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__and4_1 _3553_ (.A(_1849_),
    .B(_1852_),
    .C(_1855_),
    .D(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__and3_1 _3554_ (.A(\output_c[2][29] ),
    .B(\output_c[2][28] ),
    .C(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__xor2_1 _3555_ (.A(net80),
    .B(_1867_),
    .X(_0680_));
 sky130_fd_sc_hd__a21oi_1 _3556_ (.A1(net345),
    .A2(_1866_),
    .B1(net430),
    .Y(_1868_));
 sky130_fd_sc_hd__nor2_1 _3557_ (.A(_1867_),
    .B(_1868_),
    .Y(_0679_));
 sky130_fd_sc_hd__xor2_1 _3558_ (.A(net345),
    .B(_1866_),
    .X(_0678_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3559_ (.A(\output_c[2][24] ),
    .X(_1869_));
 sky130_fd_sc_hd__and3_1 _3560_ (.A(_1852_),
    .B(_1855_),
    .C(_1865_),
    .X(_1870_));
 sky130_fd_sc_hd__a41o_1 _3561_ (.A1(\output_c[2][26] ),
    .A2(\output_c[2][25] ),
    .A3(_1869_),
    .A4(_1870_),
    .B1(\output_c[2][27] ),
    .X(_1871_));
 sky130_fd_sc_hd__and2b_1 _3562_ (.A_N(_1866_),
    .B(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__clkbuf_1 _3563_ (.A(_1872_),
    .X(_0677_));
 sky130_fd_sc_hd__buf_1 _3564_ (.A(_1870_),
    .X(_1873_));
 sky130_fd_sc_hd__nand3_1 _3565_ (.A(\output_c[2][25] ),
    .B(_1869_),
    .C(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__xnor2_1 _3566_ (.A(net248),
    .B(_1874_),
    .Y(_0676_));
 sky130_fd_sc_hd__a21o_1 _3567_ (.A1(_1869_),
    .A2(_1873_),
    .B1(\output_c[2][25] ),
    .X(_1875_));
 sky130_fd_sc_hd__and2_1 _3568_ (.A(_1874_),
    .B(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__clkbuf_1 _3569_ (.A(_1876_),
    .X(_0675_));
 sky130_fd_sc_hd__xor2_1 _3570_ (.A(_1869_),
    .B(_1873_),
    .X(_0674_));
 sky130_fd_sc_hd__buf_1 _3571_ (.A(_1855_),
    .X(_1877_));
 sky130_fd_sc_hd__a41o_1 _3572_ (.A1(\output_c[2][22] ),
    .A2(_1851_),
    .A3(_1877_),
    .A4(_1861_),
    .B1(\output_c[2][23] ),
    .X(_1878_));
 sky130_fd_sc_hd__and2b_1 _3573_ (.A_N(_1873_),
    .B(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__clkbuf_1 _3574_ (.A(_1879_),
    .X(_0673_));
 sky130_fd_sc_hd__buf_1 _3575_ (.A(_1865_),
    .X(_1880_));
 sky130_fd_sc_hd__and3_1 _3576_ (.A(_1850_),
    .B(_1877_),
    .C(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__and3_1 _3577_ (.A(\output_c[2][21] ),
    .B(\output_c[2][20] ),
    .C(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__xor2_1 _3578_ (.A(net160),
    .B(_1882_),
    .X(_0672_));
 sky130_fd_sc_hd__a21oi_1 _3579_ (.A1(\output_c[2][20] ),
    .A2(_1881_),
    .B1(net284),
    .Y(_1883_));
 sky130_fd_sc_hd__nor2_1 _3580_ (.A(_1882_),
    .B(net285),
    .Y(_0671_));
 sky130_fd_sc_hd__xor2_1 _3581_ (.A(net331),
    .B(_1881_),
    .X(_0670_));
 sky130_fd_sc_hd__and3_1 _3582_ (.A(\output_c[2][16] ),
    .B(_1877_),
    .C(_1880_),
    .X(_1884_));
 sky130_fd_sc_hd__and3_1 _3583_ (.A(\output_c[2][18] ),
    .B(\output_c[2][17] ),
    .C(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__o21ba_1 _3584_ (.A1(net189),
    .A2(_1885_),
    .B1_N(_1881_),
    .X(_0669_));
 sky130_fd_sc_hd__a21oi_1 _3585_ (.A1(net356),
    .A2(_1884_),
    .B1(net372),
    .Y(_1886_));
 sky130_fd_sc_hd__nor2_1 _3586_ (.A(_1885_),
    .B(_1886_),
    .Y(_0668_));
 sky130_fd_sc_hd__xor2_1 _3587_ (.A(net356),
    .B(_1884_),
    .X(_0667_));
 sky130_fd_sc_hd__buf_1 _3588_ (.A(_1880_),
    .X(_1887_));
 sky130_fd_sc_hd__a21o_1 _3589_ (.A1(_1877_),
    .A2(_1887_),
    .B1(\output_c[2][16] ),
    .X(_1888_));
 sky130_fd_sc_hd__and2b_1 _3590_ (.A_N(_1884_),
    .B(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__clkbuf_1 _3591_ (.A(_1889_),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _3592_ (.A(\output_c[2][12] ),
    .B(_1853_),
    .C(_1861_),
    .X(_1890_));
 sky130_fd_sc_hd__and3_1 _3593_ (.A(\output_c[2][14] ),
    .B(\output_c[2][13] ),
    .C(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__xor2_1 _3594_ (.A(net57),
    .B(_1891_),
    .X(_0665_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3595_ (.A(_1887_),
    .X(_1892_));
 sky130_fd_sc_hd__a21oi_1 _3596_ (.A1(_1854_),
    .A2(_1892_),
    .B1(net277),
    .Y(_1893_));
 sky130_fd_sc_hd__nor2_1 _3597_ (.A(_1891_),
    .B(_1893_),
    .Y(_0664_));
 sky130_fd_sc_hd__nor2_1 _3598_ (.A(net310),
    .B(_1890_),
    .Y(_1894_));
 sky130_fd_sc_hd__a21oi_1 _3599_ (.A1(_1854_),
    .A2(_1892_),
    .B1(_1894_),
    .Y(_0663_));
 sky130_fd_sc_hd__and2_1 _3600_ (.A(_1853_),
    .B(_1887_),
    .X(_1895_));
 sky130_fd_sc_hd__nor2_1 _3601_ (.A(net341),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__nor2_1 _3602_ (.A(_1890_),
    .B(_1896_),
    .Y(_0662_));
 sky130_fd_sc_hd__and3_1 _3603_ (.A(\output_c[2][9] ),
    .B(\output_c[2][8] ),
    .C(_1880_),
    .X(_1897_));
 sky130_fd_sc_hd__a21oi_1 _3604_ (.A1(net119),
    .A2(_1897_),
    .B1(net124),
    .Y(_1898_));
 sky130_fd_sc_hd__nor2_1 _3605_ (.A(_1895_),
    .B(_1898_),
    .Y(_0661_));
 sky130_fd_sc_hd__xor2_1 _3606_ (.A(net119),
    .B(_1897_),
    .X(_0660_));
 sky130_fd_sc_hd__a21oi_1 _3607_ (.A1(net347),
    .A2(_1892_),
    .B1(net376),
    .Y(_1899_));
 sky130_fd_sc_hd__nor2_1 _3608_ (.A(_1897_),
    .B(_1899_),
    .Y(_0659_));
 sky130_fd_sc_hd__xor2_1 _3609_ (.A(net347),
    .B(_1892_),
    .X(_0658_));
 sky130_fd_sc_hd__buf_1 _3610_ (.A(_1859_),
    .X(_1900_));
 sky130_fd_sc_hd__and3_1 _3611_ (.A(\output_c[2][5] ),
    .B(_1856_),
    .C(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__a21o_1 _3612_ (.A1(\output_c[2][6] ),
    .A2(_1901_),
    .B1(\output_c[2][7] ),
    .X(_1902_));
 sky130_fd_sc_hd__and2b_1 _3613_ (.A_N(_1887_),
    .B(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_1 _3614_ (.A(_1903_),
    .X(_0657_));
 sky130_fd_sc_hd__xor2_1 _3615_ (.A(net357),
    .B(_1901_),
    .X(_0656_));
 sky130_fd_sc_hd__a21oi_1 _3616_ (.A1(_1856_),
    .A2(_1900_),
    .B1(net463),
    .Y(_1904_));
 sky130_fd_sc_hd__nor2_1 _3617_ (.A(_1901_),
    .B(_1904_),
    .Y(_0655_));
 sky130_fd_sc_hd__xor2_1 _3618_ (.A(_1856_),
    .B(_1900_),
    .X(_0654_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3619_ (.A(_1154_),
    .X(_1905_));
 sky130_fd_sc_hd__and3_1 _3620_ (.A(\output_c[2][1] ),
    .B(_1905_),
    .C(_1857_),
    .X(_1906_));
 sky130_fd_sc_hd__and2_1 _3621_ (.A(\output_c[2][2] ),
    .B(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__o21ba_1 _3622_ (.A1(net165),
    .A2(_1907_),
    .B1_N(_1900_),
    .X(_0653_));
 sky130_fd_sc_hd__nor2_1 _3623_ (.A(net350),
    .B(_1906_),
    .Y(_1908_));
 sky130_fd_sc_hd__nor2_1 _3624_ (.A(_1907_),
    .B(_1908_),
    .Y(_0652_));
 sky130_fd_sc_hd__a21oi_1 _3625_ (.A1(_1845_),
    .A2(_1857_),
    .B1(net377),
    .Y(_1909_));
 sky130_fd_sc_hd__nor2_1 _3626_ (.A(_1906_),
    .B(_1909_),
    .Y(_0651_));
 sky130_fd_sc_hd__buf_1 _3627_ (.A(_1147_),
    .X(_1910_));
 sky130_fd_sc_hd__buf_1 _3628_ (.A(_1155_),
    .X(_1911_));
 sky130_fd_sc_hd__and3_1 _3629_ (.A(_1847_),
    .B(\input_a[2][0] ),
    .C(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__o2bb2a_1 _3630_ (.A1_N(_1910_),
    .A2_N(_1857_),
    .B1(_1912_),
    .B2(net184),
    .X(_0650_));
 sky130_fd_sc_hd__and2_1 _3631_ (.A(\output_c[1][25] ),
    .B(\output_c[1][24] ),
    .X(_1913_));
 sky130_fd_sc_hd__and3_1 _3632_ (.A(\output_c[1][27] ),
    .B(\output_c[1][26] ),
    .C(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__and4_1 _3633_ (.A(\output_c[1][19] ),
    .B(\output_c[1][18] ),
    .C(\output_c[1][17] ),
    .D(\output_c[1][16] ),
    .X(_1915_));
 sky130_fd_sc_hd__and3_1 _3634_ (.A(\output_c[1][21] ),
    .B(\output_c[1][20] ),
    .C(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__and3_1 _3635_ (.A(\output_c[1][23] ),
    .B(\output_c[1][22] ),
    .C(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__and4_1 _3636_ (.A(\output_c[1][11] ),
    .B(\output_c[1][10] ),
    .C(\output_c[1][9] ),
    .D(\output_c[1][8] ),
    .X(_1918_));
 sky130_fd_sc_hd__and3_1 _3637_ (.A(\output_c[1][15] ),
    .B(\output_c[1][14] ),
    .C(\output_c[1][13] ),
    .X(_1919_));
 sky130_fd_sc_hd__and3_1 _3638_ (.A(\output_c[1][12] ),
    .B(_1918_),
    .C(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__buf_1 _3639_ (.A(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__and3_1 _3640_ (.A(\output_c[1][0] ),
    .B(_1487_),
    .C(\input_a[1][0] ),
    .X(_1922_));
 sky130_fd_sc_hd__and2_1 _3641_ (.A(\output_c[1][3] ),
    .B(\output_c[1][2] ),
    .X(_1923_));
 sky130_fd_sc_hd__and4_1 _3642_ (.A(\output_c[1][1] ),
    .B(_1101_),
    .C(_1922_),
    .D(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__and2_1 _3643_ (.A(\output_c[1][7] ),
    .B(\output_c[1][6] ),
    .X(_1925_));
 sky130_fd_sc_hd__and4_1 _3644_ (.A(\output_c[1][5] ),
    .B(\output_c[1][4] ),
    .C(_1924_),
    .D(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__and4_1 _3645_ (.A(_1914_),
    .B(_1917_),
    .C(_1921_),
    .D(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__and4_1 _3646_ (.A(\output_c[1][30] ),
    .B(\output_c[1][29] ),
    .C(\output_c[1][28] ),
    .D(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__xor2_1 _3647_ (.A(net36),
    .B(_1928_),
    .X(_0649_));
 sky130_fd_sc_hd__buf_1 _3648_ (.A(\output_c[1][4] ),
    .X(_1929_));
 sky130_fd_sc_hd__and2_1 _3649_ (.A(\output_c[1][6] ),
    .B(\output_c[1][5] ),
    .X(_1930_));
 sky130_fd_sc_hd__and4_1 _3650_ (.A(\output_c[1][7] ),
    .B(_1929_),
    .C(_1924_),
    .D(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__and4_2 _3651_ (.A(_1914_),
    .B(_1917_),
    .C(_1920_),
    .D(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__and3_1 _3652_ (.A(\output_c[1][29] ),
    .B(\output_c[1][28] ),
    .C(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__xor2_1 _3653_ (.A(net59),
    .B(_1933_),
    .X(_0648_));
 sky130_fd_sc_hd__a21oi_1 _3654_ (.A1(\output_c[1][28] ),
    .A2(_1932_),
    .B1(net342),
    .Y(_1934_));
 sky130_fd_sc_hd__nor2_1 _3655_ (.A(_1933_),
    .B(net343),
    .Y(_0647_));
 sky130_fd_sc_hd__xor2_1 _3656_ (.A(net359),
    .B(_1932_),
    .X(_0646_));
 sky130_fd_sc_hd__buf_1 _3657_ (.A(_1917_),
    .X(_1935_));
 sky130_fd_sc_hd__buf_1 _3658_ (.A(_1931_),
    .X(_1936_));
 sky130_fd_sc_hd__and4_1 _3659_ (.A(_1913_),
    .B(_1935_),
    .C(_1921_),
    .D(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__a21oi_1 _3660_ (.A1(\output_c[1][26] ),
    .A2(_1937_),
    .B1(net117),
    .Y(_1938_));
 sky130_fd_sc_hd__nor2_1 _3661_ (.A(_1932_),
    .B(net118),
    .Y(_0645_));
 sky130_fd_sc_hd__xor2_1 _3662_ (.A(net162),
    .B(_1937_),
    .X(_0644_));
 sky130_fd_sc_hd__and2_1 _3663_ (.A(_1920_),
    .B(_1926_),
    .X(_1939_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3664_ (.A(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__nand3_1 _3665_ (.A(\output_c[1][24] ),
    .B(_1935_),
    .C(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__xnor2_1 _3666_ (.A(net74),
    .B(_1941_),
    .Y(_0643_));
 sky130_fd_sc_hd__a31o_1 _3667_ (.A1(_1935_),
    .A2(_1921_),
    .A3(_1936_),
    .B1(\output_c[1][24] ),
    .X(_1942_));
 sky130_fd_sc_hd__and2_1 _3668_ (.A(_1941_),
    .B(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__clkbuf_1 _3669_ (.A(_1943_),
    .X(_0642_));
 sky130_fd_sc_hd__a31o_1 _3670_ (.A1(\output_c[1][22] ),
    .A2(_1916_),
    .A3(_1940_),
    .B1(net486),
    .X(_1944_));
 sky130_fd_sc_hd__a21boi_1 _3671_ (.A1(_1935_),
    .A2(_1940_),
    .B1_N(net487),
    .Y(_0641_));
 sky130_fd_sc_hd__and3_1 _3672_ (.A(_1915_),
    .B(_1921_),
    .C(_1931_),
    .X(_1945_));
 sky130_fd_sc_hd__and3_1 _3673_ (.A(\output_c[1][21] ),
    .B(\output_c[1][20] ),
    .C(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__xor2_1 _3674_ (.A(net101),
    .B(_1946_),
    .X(_0640_));
 sky130_fd_sc_hd__a21oi_1 _3675_ (.A1(\output_c[1][20] ),
    .A2(_1945_),
    .B1(net221),
    .Y(_1947_));
 sky130_fd_sc_hd__nor2_1 _3676_ (.A(_1946_),
    .B(net222),
    .Y(_0639_));
 sky130_fd_sc_hd__xor2_1 _3677_ (.A(net266),
    .B(_1945_),
    .X(_0638_));
 sky130_fd_sc_hd__and3_1 _3678_ (.A(\output_c[1][16] ),
    .B(_1920_),
    .C(_1931_),
    .X(_1948_));
 sky130_fd_sc_hd__a31o_1 _3679_ (.A1(\output_c[1][18] ),
    .A2(\output_c[1][17] ),
    .A3(_1948_),
    .B1(\output_c[1][19] ),
    .X(_1949_));
 sky130_fd_sc_hd__and2b_1 _3680_ (.A_N(_1945_),
    .B(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__clkbuf_1 _3681_ (.A(_1950_),
    .X(_0637_));
 sky130_fd_sc_hd__and3_1 _3682_ (.A(\output_c[1][17] ),
    .B(\output_c[1][16] ),
    .C(_1939_),
    .X(_1951_));
 sky130_fd_sc_hd__xor2_1 _3683_ (.A(net171),
    .B(_1951_),
    .X(_0636_));
 sky130_fd_sc_hd__nor2_1 _3684_ (.A(net481),
    .B(_1948_),
    .Y(_1952_));
 sky130_fd_sc_hd__nor2_1 _3685_ (.A(_1951_),
    .B(_1952_),
    .Y(_0635_));
 sky130_fd_sc_hd__xor2_1 _3686_ (.A(net217),
    .B(_1940_),
    .X(_0634_));
 sky130_fd_sc_hd__and3_1 _3687_ (.A(\output_c[1][12] ),
    .B(_1918_),
    .C(_1926_),
    .X(_1953_));
 sky130_fd_sc_hd__and3_1 _3688_ (.A(\output_c[1][14] ),
    .B(\output_c[1][13] ),
    .C(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__xor2_1 _3689_ (.A(net79),
    .B(_1954_),
    .X(_0633_));
 sky130_fd_sc_hd__a21o_1 _3690_ (.A1(\output_c[1][13] ),
    .A2(_1953_),
    .B1(\output_c[1][14] ),
    .X(_1955_));
 sky130_fd_sc_hd__and2b_1 _3691_ (.A_N(_1954_),
    .B(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__clkbuf_1 _3692_ (.A(_1956_),
    .X(_0632_));
 sky130_fd_sc_hd__xor2_1 _3693_ (.A(net407),
    .B(_1953_),
    .X(_0631_));
 sky130_fd_sc_hd__buf_1 _3694_ (.A(_1936_),
    .X(_1957_));
 sky130_fd_sc_hd__and2_1 _3695_ (.A(_1918_),
    .B(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__nor2_1 _3696_ (.A(net433),
    .B(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nor2_1 _3697_ (.A(_1953_),
    .B(_1959_),
    .Y(_0630_));
 sky130_fd_sc_hd__and3_1 _3698_ (.A(\output_c[1][9] ),
    .B(\output_c[1][8] ),
    .C(_1936_),
    .X(_1960_));
 sky130_fd_sc_hd__a21oi_1 _3699_ (.A1(net212),
    .A2(_1960_),
    .B1(net219),
    .Y(_1961_));
 sky130_fd_sc_hd__nor2_1 _3700_ (.A(_1958_),
    .B(_1961_),
    .Y(_0629_));
 sky130_fd_sc_hd__xor2_1 _3701_ (.A(net212),
    .B(_1960_),
    .X(_0628_));
 sky130_fd_sc_hd__a21oi_1 _3702_ (.A1(net378),
    .A2(_1957_),
    .B1(net403),
    .Y(_1962_));
 sky130_fd_sc_hd__nor2_1 _3703_ (.A(_1960_),
    .B(_1962_),
    .Y(_0627_));
 sky130_fd_sc_hd__xor2_1 _3704_ (.A(net378),
    .B(_1957_),
    .X(_0626_));
 sky130_fd_sc_hd__buf_1 _3705_ (.A(_1924_),
    .X(_1963_));
 sky130_fd_sc_hd__and3_1 _3706_ (.A(\output_c[1][5] ),
    .B(_1929_),
    .C(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__a21o_1 _3707_ (.A1(\output_c[1][6] ),
    .A2(_1964_),
    .B1(\output_c[1][7] ),
    .X(_1965_));
 sky130_fd_sc_hd__and2b_1 _3708_ (.A_N(_1957_),
    .B(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__clkbuf_1 _3709_ (.A(_1966_),
    .X(_0625_));
 sky130_fd_sc_hd__xor2_1 _3710_ (.A(net262),
    .B(_1964_),
    .X(_0624_));
 sky130_fd_sc_hd__a21oi_1 _3711_ (.A1(_1929_),
    .A2(_1963_),
    .B1(net475),
    .Y(_1967_));
 sky130_fd_sc_hd__nor2_1 _3712_ (.A(_1964_),
    .B(_1967_),
    .Y(_0623_));
 sky130_fd_sc_hd__xor2_1 _3713_ (.A(_1929_),
    .B(_1963_),
    .X(_0622_));
 sky130_fd_sc_hd__and3_1 _3714_ (.A(\output_c[1][1] ),
    .B(_1905_),
    .C(_1922_),
    .X(_1968_));
 sky130_fd_sc_hd__and2_1 _3715_ (.A(\output_c[1][2] ),
    .B(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__o21ba_1 _3716_ (.A1(net169),
    .A2(_1969_),
    .B1_N(_1963_),
    .X(_0621_));
 sky130_fd_sc_hd__nor2_1 _3717_ (.A(net442),
    .B(_1968_),
    .Y(_1970_));
 sky130_fd_sc_hd__nor2_1 _3718_ (.A(_1969_),
    .B(_1970_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21oi_1 _3719_ (.A1(_1845_),
    .A2(_1922_),
    .B1(net375),
    .Y(_1971_));
 sky130_fd_sc_hd__nor2_1 _3720_ (.A(_1968_),
    .B(_1971_),
    .Y(_0619_));
 sky130_fd_sc_hd__and3_1 _3721_ (.A(_1847_),
    .B(\input_a[1][0] ),
    .C(_1911_),
    .X(_1972_));
 sky130_fd_sc_hd__o2bb2a_1 _3722_ (.A1_N(_1910_),
    .A2_N(_1922_),
    .B1(_1972_),
    .B2(net167),
    .X(_0618_));
 sky130_fd_sc_hd__and4_1 _3723_ (.A(\output_c[0][27] ),
    .B(\output_c[0][26] ),
    .C(\output_c[0][25] ),
    .D(\output_c[0][24] ),
    .X(_1973_));
 sky130_fd_sc_hd__and4_1 _3724_ (.A(\output_c[0][19] ),
    .B(\output_c[0][18] ),
    .C(\output_c[0][17] ),
    .D(\output_c[0][16] ),
    .X(_1974_));
 sky130_fd_sc_hd__and3_1 _3725_ (.A(\output_c[0][21] ),
    .B(\output_c[0][20] ),
    .C(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__and3_1 _3726_ (.A(\output_c[0][23] ),
    .B(\output_c[0][22] ),
    .C(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__buf_1 _3727_ (.A(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__and4_1 _3728_ (.A(\output_c[0][11] ),
    .B(\output_c[0][10] ),
    .C(\output_c[0][9] ),
    .D(\output_c[0][8] ),
    .X(_1978_));
 sky130_fd_sc_hd__and3_1 _3729_ (.A(\output_c[0][13] ),
    .B(\output_c[0][12] ),
    .C(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__and3_1 _3730_ (.A(\output_c[0][15] ),
    .B(\output_c[0][14] ),
    .C(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__buf_1 _3731_ (.A(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__buf_1 _3732_ (.A(\output_c[0][4] ),
    .X(_1982_));
 sky130_fd_sc_hd__and3_1 _3733_ (.A(\output_c[0][0] ),
    .B(_1289_),
    .C(\input_a[0][0] ),
    .X(_1983_));
 sky130_fd_sc_hd__and2_1 _3734_ (.A(\output_c[0][3] ),
    .B(\output_c[0][2] ),
    .X(_1984_));
 sky130_fd_sc_hd__and4_1 _3735_ (.A(\output_c[0][1] ),
    .B(_1164_),
    .C(_1983_),
    .D(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__and2_1 _3736_ (.A(\output_c[0][7] ),
    .B(\output_c[0][6] ),
    .X(_1986_));
 sky130_fd_sc_hd__and4_1 _3737_ (.A(\output_c[0][5] ),
    .B(_1982_),
    .C(_1985_),
    .D(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__and4_1 _3738_ (.A(_1973_),
    .B(_1977_),
    .C(_1981_),
    .D(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__and4_1 _3739_ (.A(\output_c[0][30] ),
    .B(\output_c[0][29] ),
    .C(\output_c[0][28] ),
    .D(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__xor2_1 _3740_ (.A(net48),
    .B(_1989_),
    .X(_0617_));
 sky130_fd_sc_hd__and2_1 _3741_ (.A(\output_c[0][6] ),
    .B(\output_c[0][5] ),
    .X(_1990_));
 sky130_fd_sc_hd__and4_1 _3742_ (.A(\output_c[0][7] ),
    .B(\output_c[0][4] ),
    .C(_1985_),
    .D(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__buf_1 _3743_ (.A(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__and4_1 _3744_ (.A(_1973_),
    .B(_1977_),
    .C(_1981_),
    .D(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__and3_1 _3745_ (.A(\output_c[0][29] ),
    .B(\output_c[0][28] ),
    .C(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__xor2_1 _3746_ (.A(net90),
    .B(_1994_),
    .X(_0616_));
 sky130_fd_sc_hd__a21oi_1 _3747_ (.A1(net390),
    .A2(_1993_),
    .B1(net435),
    .Y(_1995_));
 sky130_fd_sc_hd__nor2_1 _3748_ (.A(_1994_),
    .B(_1995_),
    .Y(_0615_));
 sky130_fd_sc_hd__xor2_1 _3749_ (.A(net390),
    .B(_1993_),
    .X(_0614_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3750_ (.A(\output_c[0][24] ),
    .X(_1996_));
 sky130_fd_sc_hd__and3_1 _3751_ (.A(_1976_),
    .B(_1980_),
    .C(_1991_),
    .X(_1997_));
 sky130_fd_sc_hd__a41o_1 _3752_ (.A1(\output_c[0][26] ),
    .A2(\output_c[0][25] ),
    .A3(_1996_),
    .A4(_1997_),
    .B1(\output_c[0][27] ),
    .X(_1998_));
 sky130_fd_sc_hd__and2b_1 _3753_ (.A_N(_1993_),
    .B(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__clkbuf_1 _3754_ (.A(_1999_),
    .X(_0613_));
 sky130_fd_sc_hd__and2_1 _3755_ (.A(_1980_),
    .B(_1987_),
    .X(_2000_));
 sky130_fd_sc_hd__and4_1 _3756_ (.A(\output_c[0][25] ),
    .B(_1996_),
    .C(_1977_),
    .D(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__xor2_1 _3757_ (.A(net329),
    .B(_2001_),
    .X(_0612_));
 sky130_fd_sc_hd__a21o_1 _3758_ (.A1(_1996_),
    .A2(_1997_),
    .B1(\output_c[0][25] ),
    .X(_2002_));
 sky130_fd_sc_hd__and2b_1 _3759_ (.A_N(_2001_),
    .B(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__clkbuf_1 _3760_ (.A(_2003_),
    .X(_0611_));
 sky130_fd_sc_hd__xor2_1 _3761_ (.A(_1996_),
    .B(_1997_),
    .X(_0610_));
 sky130_fd_sc_hd__buf_1 _3762_ (.A(_2000_),
    .X(_2004_));
 sky130_fd_sc_hd__a31o_1 _3763_ (.A1(\output_c[0][22] ),
    .A2(_1975_),
    .A3(_2004_),
    .B1(net489),
    .X(_2005_));
 sky130_fd_sc_hd__a21boi_1 _3764_ (.A1(_1977_),
    .A2(_2004_),
    .B1_N(_2005_),
    .Y(_0609_));
 sky130_fd_sc_hd__and3_1 _3765_ (.A(_1974_),
    .B(_1981_),
    .C(_1992_),
    .X(_2006_));
 sky130_fd_sc_hd__and3_1 _3766_ (.A(\output_c[0][21] ),
    .B(\output_c[0][20] ),
    .C(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__xor2_1 _3767_ (.A(net96),
    .B(_2007_),
    .X(_0608_));
 sky130_fd_sc_hd__a21oi_1 _3768_ (.A1(net327),
    .A2(_2006_),
    .B1(net361),
    .Y(_2008_));
 sky130_fd_sc_hd__nor2_1 _3769_ (.A(_2007_),
    .B(_2008_),
    .Y(_0607_));
 sky130_fd_sc_hd__xor2_1 _3770_ (.A(net327),
    .B(_2006_),
    .X(_0606_));
 sky130_fd_sc_hd__and3_1 _3771_ (.A(\output_c[0][16] ),
    .B(_1981_),
    .C(_1992_),
    .X(_2009_));
 sky130_fd_sc_hd__a31o_1 _3772_ (.A1(\output_c[0][18] ),
    .A2(\output_c[0][17] ),
    .A3(_2009_),
    .B1(\output_c[0][19] ),
    .X(_2010_));
 sky130_fd_sc_hd__and2b_1 _3773_ (.A_N(_2006_),
    .B(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__clkbuf_1 _3774_ (.A(_2011_),
    .X(_0605_));
 sky130_fd_sc_hd__and3_1 _3775_ (.A(\output_c[0][17] ),
    .B(\output_c[0][16] ),
    .C(_2004_),
    .X(_2012_));
 sky130_fd_sc_hd__xor2_1 _3776_ (.A(net158),
    .B(_2012_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _3777_ (.A(net479),
    .B(_2009_),
    .Y(_2013_));
 sky130_fd_sc_hd__nor2_1 _3778_ (.A(_2012_),
    .B(_2013_),
    .Y(_0603_));
 sky130_fd_sc_hd__xor2_1 _3779_ (.A(net237),
    .B(_2004_),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _3780_ (.A(\output_c[0][12] ),
    .B(_1978_),
    .C(_1987_),
    .X(_2014_));
 sky130_fd_sc_hd__and3_1 _3781_ (.A(\output_c[0][14] ),
    .B(\output_c[0][13] ),
    .C(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__xor2_1 _3782_ (.A(net66),
    .B(_2015_),
    .X(_0601_));
 sky130_fd_sc_hd__buf_1 _3783_ (.A(_1992_),
    .X(_2016_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3784_ (.A(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__a21oi_1 _3785_ (.A1(_1979_),
    .A2(_2017_),
    .B1(net409),
    .Y(_2018_));
 sky130_fd_sc_hd__nor2_1 _3786_ (.A(_2015_),
    .B(_2018_),
    .Y(_0600_));
 sky130_fd_sc_hd__nor2_1 _3787_ (.A(net332),
    .B(_2014_),
    .Y(_2019_));
 sky130_fd_sc_hd__a21oi_1 _3788_ (.A1(_1979_),
    .A2(_2017_),
    .B1(_2019_),
    .Y(_0599_));
 sky130_fd_sc_hd__and2_1 _3789_ (.A(_1978_),
    .B(_2016_),
    .X(_2020_));
 sky130_fd_sc_hd__nor2_1 _3790_ (.A(net422),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__nor2_1 _3791_ (.A(_2014_),
    .B(_2021_),
    .Y(_0598_));
 sky130_fd_sc_hd__and3_1 _3792_ (.A(\output_c[0][9] ),
    .B(\output_c[0][8] ),
    .C(_2016_),
    .X(_2022_));
 sky130_fd_sc_hd__a21oi_1 _3793_ (.A1(net127),
    .A2(_2022_),
    .B1(net146),
    .Y(_2023_));
 sky130_fd_sc_hd__nor2_1 _3794_ (.A(_2020_),
    .B(_2023_),
    .Y(_0597_));
 sky130_fd_sc_hd__xor2_1 _3795_ (.A(net127),
    .B(_2022_),
    .X(_0596_));
 sky130_fd_sc_hd__a21oi_1 _3796_ (.A1(net298),
    .A2(_2017_),
    .B1(net416),
    .Y(_2024_));
 sky130_fd_sc_hd__nor2_1 _3797_ (.A(_2022_),
    .B(_2024_),
    .Y(_0595_));
 sky130_fd_sc_hd__xor2_1 _3798_ (.A(net298),
    .B(_2017_),
    .X(_0594_));
 sky130_fd_sc_hd__buf_1 _3799_ (.A(_1985_),
    .X(_2025_));
 sky130_fd_sc_hd__and3_1 _3800_ (.A(\output_c[0][5] ),
    .B(_1982_),
    .C(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__a21o_1 _3801_ (.A1(\output_c[0][6] ),
    .A2(_2026_),
    .B1(\output_c[0][7] ),
    .X(_2027_));
 sky130_fd_sc_hd__and2b_1 _3802_ (.A_N(_2016_),
    .B(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__clkbuf_1 _3803_ (.A(_2028_),
    .X(_0593_));
 sky130_fd_sc_hd__xor2_1 _3804_ (.A(net379),
    .B(_2026_),
    .X(_0592_));
 sky130_fd_sc_hd__a21oi_1 _3805_ (.A1(_1982_),
    .A2(_2025_),
    .B1(net473),
    .Y(_2029_));
 sky130_fd_sc_hd__nor2_1 _3806_ (.A(_2026_),
    .B(_2029_),
    .Y(_0591_));
 sky130_fd_sc_hd__xor2_1 _3807_ (.A(_1982_),
    .B(_2025_),
    .X(_0590_));
 sky130_fd_sc_hd__and3_1 _3808_ (.A(\output_c[0][1] ),
    .B(_1905_),
    .C(_1983_),
    .X(_2030_));
 sky130_fd_sc_hd__and2_1 _3809_ (.A(\output_c[0][2] ),
    .B(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__o21ba_1 _3810_ (.A1(net200),
    .A2(_2031_),
    .B1_N(_2025_),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _3811_ (.A(net413),
    .B(_2030_),
    .Y(_2032_));
 sky130_fd_sc_hd__nor2_1 _3812_ (.A(_2031_),
    .B(_2032_),
    .Y(_0588_));
 sky130_fd_sc_hd__a21oi_1 _3813_ (.A1(_1845_),
    .A2(_1983_),
    .B1(net393),
    .Y(_2033_));
 sky130_fd_sc_hd__nor2_1 _3814_ (.A(_2030_),
    .B(_2033_),
    .Y(_0587_));
 sky130_fd_sc_hd__and3_1 _3815_ (.A(_1847_),
    .B(\input_a[0][0] ),
    .C(_1911_),
    .X(_2034_));
 sky130_fd_sc_hd__o2bb2a_1 _3816_ (.A1_N(_1910_),
    .A2_N(_1983_),
    .B1(_2034_),
    .B2(net177),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_1 _3817_ (.A(_1153_),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _3818_ (.A(_2035_),
    .X(_0585_));
 sky130_fd_sc_hd__buf_1 _3819_ (.A(net1),
    .X(_2036_));
 sky130_fd_sc_hd__buf_1 _3820_ (.A(\state[2] ),
    .X(_2037_));
 sky130_fd_sc_hd__buf_1 _3821_ (.A(\state[3] ),
    .X(_2038_));
 sky130_fd_sc_hd__nand2_1 _3822_ (.A(_2037_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__buf_1 _3823_ (.A(\state[1] ),
    .X(_2040_));
 sky130_fd_sc_hd__inv_2 _3824_ (.A(net60),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2_1 _3825_ (.A(_2040_),
    .B(_0000_),
    .Y(_2041_));
 sky130_fd_sc_hd__buf_1 _3826_ (.A(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__nor2_1 _3827_ (.A(_2039_),
    .B(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__mux2_1 _3828_ (.A0(\input_a[13][0] ),
    .A1(_2036_),
    .S(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _3829_ (.A(_2044_),
    .X(_0584_));
 sky130_fd_sc_hd__or2_1 _3830_ (.A(_2040_),
    .B(_0000_),
    .X(_2045_));
 sky130_fd_sc_hd__nor2_1 _3831_ (.A(_2039_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(\input_a[12][0] ),
    .A1(_2036_),
    .S(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__clkbuf_1 _3833_ (.A(_2047_),
    .X(_0583_));
 sky130_fd_sc_hd__buf_1 _3834_ (.A(net1),
    .X(_2048_));
 sky130_fd_sc_hd__buf_1 _3835_ (.A(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__buf_1 _3836_ (.A(_2040_),
    .X(_2050_));
 sky130_fd_sc_hd__buf_1 _3837_ (.A(\state[0] ),
    .X(_2051_));
 sky130_fd_sc_hd__buf_1 _3838_ (.A(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__or3_1 _3839_ (.A(_2050_),
    .B(_2052_),
    .C(_2039_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2_1 _3840_ (.A0(_2049_),
    .A1(\input_a[11][0] ),
    .S(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _3841_ (.A(_2054_),
    .X(_0582_));
 sky130_fd_sc_hd__buf_1 _3842_ (.A(_2037_),
    .X(_2055_));
 sky130_fd_sc_hd__buf_1 _3843_ (.A(_2038_),
    .X(_2056_));
 sky130_fd_sc_hd__and4b_1 _3844_ (.A_N(_2055_),
    .B(_2056_),
    .C(_2050_),
    .D(_2052_),
    .X(_2057_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(\input_a[10][0] ),
    .A1(_2048_),
    .S(_2057_),
    .X(_2058_));
 sky130_fd_sc_hd__clkbuf_1 _3846_ (.A(_2058_),
    .X(_0581_));
 sky130_fd_sc_hd__buf_1 _3847_ (.A(_2037_),
    .X(_2059_));
 sky130_fd_sc_hd__buf_1 _3848_ (.A(_2038_),
    .X(_2060_));
 sky130_fd_sc_hd__or3b_1 _3849_ (.A(_2041_),
    .B(_2059_),
    .C_N(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__mux2_1 _3850_ (.A0(_2049_),
    .A1(\input_a[9][0] ),
    .S(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _3851_ (.A(_2062_),
    .X(_0580_));
 sky130_fd_sc_hd__or3b_1 _3852_ (.A(_2045_),
    .B(_2059_),
    .C_N(_2060_),
    .X(_2063_));
 sky130_fd_sc_hd__mux2_1 _3853_ (.A0(_2049_),
    .A1(\input_a[8][0] ),
    .S(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _3854_ (.A(_2064_),
    .X(_0579_));
 sky130_fd_sc_hd__buf_1 _3855_ (.A(_2040_),
    .X(_2065_));
 sky130_fd_sc_hd__buf_1 _3856_ (.A(_2038_),
    .X(_2066_));
 sky130_fd_sc_hd__or4b_1 _3857_ (.A(_2065_),
    .B(_2051_),
    .C(_2037_),
    .D_N(_2066_),
    .X(_2067_));
 sky130_fd_sc_hd__mux2_1 _3858_ (.A0(_2049_),
    .A1(\input_a[7][0] ),
    .S(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__clkbuf_1 _3859_ (.A(_2068_),
    .X(_0578_));
 sky130_fd_sc_hd__and4b_1 _3860_ (.A_N(_2056_),
    .B(_2055_),
    .C(_2052_),
    .D(_2050_),
    .X(_2069_));
 sky130_fd_sc_hd__mux2_1 _3861_ (.A0(\input_a[6][0] ),
    .A1(_2048_),
    .S(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__clkbuf_1 _3862_ (.A(_2070_),
    .X(_0577_));
 sky130_fd_sc_hd__buf_1 _3863_ (.A(net1),
    .X(_2071_));
 sky130_fd_sc_hd__or3b_1 _3864_ (.A(_2060_),
    .B(_2042_),
    .C_N(_2059_),
    .X(_2072_));
 sky130_fd_sc_hd__mux2_1 _3865_ (.A0(_2071_),
    .A1(\input_a[5][0] ),
    .S(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__clkbuf_1 _3866_ (.A(_2073_),
    .X(_0576_));
 sky130_fd_sc_hd__or3b_1 _3867_ (.A(_2060_),
    .B(_2045_),
    .C_N(_2059_),
    .X(_2074_));
 sky130_fd_sc_hd__mux2_1 _3868_ (.A0(_2071_),
    .A1(\input_a[4][0] ),
    .S(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__clkbuf_1 _3869_ (.A(_2075_),
    .X(_0575_));
 sky130_fd_sc_hd__buf_1 _3870_ (.A(\state[2] ),
    .X(_2076_));
 sky130_fd_sc_hd__or4b_1 _3871_ (.A(_2065_),
    .B(_2051_),
    .C(_2066_),
    .D_N(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__mux2_1 _3872_ (.A0(_2071_),
    .A1(\input_a[3][0] ),
    .S(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__clkbuf_1 _3873_ (.A(_2078_),
    .X(_0574_));
 sky130_fd_sc_hd__nand2_1 _3874_ (.A(_2065_),
    .B(_2051_),
    .Y(_2079_));
 sky130_fd_sc_hd__or3_1 _3875_ (.A(_2076_),
    .B(_2066_),
    .C(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(_2071_),
    .A1(\input_a[2][0] ),
    .S(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__clkbuf_1 _3877_ (.A(_2081_),
    .X(_0573_));
 sky130_fd_sc_hd__or3_1 _3878_ (.A(_2076_),
    .B(_2066_),
    .C(_2042_),
    .X(_2082_));
 sky130_fd_sc_hd__mux2_1 _3879_ (.A0(_2036_),
    .A1(\input_a[1][0] ),
    .S(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__clkbuf_1 _3880_ (.A(_2083_),
    .X(_0572_));
 sky130_fd_sc_hd__or3_1 _3881_ (.A(_2065_),
    .B(_2076_),
    .C(_2056_),
    .X(_2084_));
 sky130_fd_sc_hd__mux2_1 _3882_ (.A0(_2036_),
    .A1(\input_a[0][0] ),
    .S(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__clkbuf_1 _3883_ (.A(_2085_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _3884_ (.A(net490),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_1 _3885_ (.A(_2086_),
    .X(_0570_));
 sky130_fd_sc_hd__and4_1 _3886_ (.A(\output_c[15][27] ),
    .B(\output_c[15][26] ),
    .C(\output_c[15][25] ),
    .D(\output_c[15][24] ),
    .X(_2087_));
 sky130_fd_sc_hd__and4_1 _3887_ (.A(\output_c[15][19] ),
    .B(\output_c[15][18] ),
    .C(\output_c[15][17] ),
    .D(\output_c[15][16] ),
    .X(_2088_));
 sky130_fd_sc_hd__and3_1 _3888_ (.A(\output_c[15][21] ),
    .B(\output_c[15][20] ),
    .C(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__and3_1 _3889_ (.A(\output_c[15][23] ),
    .B(\output_c[15][22] ),
    .C(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__and3_1 _3890_ (.A(_1487_),
    .B(\input_a[15] ),
    .C(\output_c[15][0] ),
    .X(_2091_));
 sky130_fd_sc_hd__and2_1 _3891_ (.A(\output_c[15][3] ),
    .B(\output_c[15][2] ),
    .X(_2092_));
 sky130_fd_sc_hd__and4_1 _3892_ (.A(\output_c[15][1] ),
    .B(_1079_),
    .C(_2091_),
    .D(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__and2_1 _3893_ (.A(\output_c[15][7] ),
    .B(\output_c[15][6] ),
    .X(_2094_));
 sky130_fd_sc_hd__and4_1 _3894_ (.A(\output_c[15][5] ),
    .B(\output_c[15][4] ),
    .C(_2093_),
    .D(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__buf_1 _3895_ (.A(_2095_),
    .X(_2096_));
 sky130_fd_sc_hd__and4_1 _3896_ (.A(\output_c[15][11] ),
    .B(\output_c[15][10] ),
    .C(\output_c[15][9] ),
    .D(\output_c[15][8] ),
    .X(_2097_));
 sky130_fd_sc_hd__and3_1 _3897_ (.A(\output_c[15][13] ),
    .B(\output_c[15][12] ),
    .C(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__and3_1 _3898_ (.A(\output_c[15][15] ),
    .B(\output_c[15][14] ),
    .C(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__buf_1 _3899_ (.A(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__and4_1 _3900_ (.A(_2087_),
    .B(_2090_),
    .C(_2096_),
    .D(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__and4_1 _3901_ (.A(\output_c[15][30] ),
    .B(\output_c[15][29] ),
    .C(\output_c[15][28] ),
    .D(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__xor2_1 _3902_ (.A(net50),
    .B(_2102_),
    .X(_0569_));
 sky130_fd_sc_hd__buf_1 _3903_ (.A(\output_c[15][4] ),
    .X(_2103_));
 sky130_fd_sc_hd__and2_1 _3904_ (.A(\output_c[15][6] ),
    .B(\output_c[15][5] ),
    .X(_2104_));
 sky130_fd_sc_hd__and4_1 _3905_ (.A(\output_c[15][7] ),
    .B(_2103_),
    .C(_2093_),
    .D(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__and4_1 _3906_ (.A(_2087_),
    .B(_2090_),
    .C(_2100_),
    .D(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__and3_1 _3907_ (.A(\output_c[15][29] ),
    .B(\output_c[15][28] ),
    .C(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__xor2_1 _3908_ (.A(net77),
    .B(_2107_),
    .X(_0568_));
 sky130_fd_sc_hd__a21oi_1 _3909_ (.A1(net338),
    .A2(_2106_),
    .B1(net400),
    .Y(_2108_));
 sky130_fd_sc_hd__nor2_1 _3910_ (.A(_2107_),
    .B(_2108_),
    .Y(_0567_));
 sky130_fd_sc_hd__xor2_1 _3911_ (.A(net338),
    .B(_2106_),
    .X(_0566_));
 sky130_fd_sc_hd__and4_1 _3912_ (.A(\output_c[15][24] ),
    .B(_2090_),
    .C(_2096_),
    .D(_2100_),
    .X(_2109_));
 sky130_fd_sc_hd__and3_1 _3913_ (.A(\output_c[15][26] ),
    .B(\output_c[15][25] ),
    .C(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__o21ba_1 _3914_ (.A1(net257),
    .A2(_2110_),
    .B1_N(_2106_),
    .X(_0565_));
 sky130_fd_sc_hd__nand2_1 _3915_ (.A(net494),
    .B(_2109_),
    .Y(_2111_));
 sky130_fd_sc_hd__xnor2_1 _3916_ (.A(net175),
    .B(_2111_),
    .Y(_0564_));
 sky130_fd_sc_hd__xor2_1 _3917_ (.A(net307),
    .B(_2109_),
    .X(_0563_));
 sky130_fd_sc_hd__buf_1 _3918_ (.A(_2100_),
    .X(_2112_));
 sky130_fd_sc_hd__buf_1 _3919_ (.A(_2105_),
    .X(_2113_));
 sky130_fd_sc_hd__a31o_1 _3920_ (.A1(_2090_),
    .A2(_2112_),
    .A3(_2113_),
    .B1(\output_c[15][24] ),
    .X(_2114_));
 sky130_fd_sc_hd__and2b_1 _3921_ (.A_N(_2109_),
    .B(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__clkbuf_1 _3922_ (.A(_2115_),
    .X(_0562_));
 sky130_fd_sc_hd__and4_1 _3923_ (.A(\output_c[15][22] ),
    .B(_2089_),
    .C(_2096_),
    .D(_2112_),
    .X(_2116_));
 sky130_fd_sc_hd__xor2_1 _3924_ (.A(net67),
    .B(_2116_),
    .X(_0561_));
 sky130_fd_sc_hd__and3_1 _3925_ (.A(_2088_),
    .B(_2099_),
    .C(_2105_),
    .X(_2117_));
 sky130_fd_sc_hd__nand3_1 _3926_ (.A(\output_c[15][21] ),
    .B(\output_c[15][20] ),
    .C(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__xnor2_1 _3927_ (.A(net144),
    .B(_2118_),
    .Y(_0560_));
 sky130_fd_sc_hd__a21o_1 _3928_ (.A1(\output_c[15][20] ),
    .A2(_2117_),
    .B1(\output_c[15][21] ),
    .X(_2119_));
 sky130_fd_sc_hd__and2_1 _3929_ (.A(_2118_),
    .B(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__clkbuf_1 _3930_ (.A(_2120_),
    .X(_0559_));
 sky130_fd_sc_hd__xor2_1 _3931_ (.A(net426),
    .B(_2117_),
    .X(_0558_));
 sky130_fd_sc_hd__and4_1 _3932_ (.A(\output_c[15][17] ),
    .B(\output_c[15][16] ),
    .C(_2095_),
    .D(_2099_),
    .X(_2121_));
 sky130_fd_sc_hd__a21o_1 _3933_ (.A1(\output_c[15][18] ),
    .A2(_2121_),
    .B1(\output_c[15][19] ),
    .X(_2122_));
 sky130_fd_sc_hd__and2b_1 _3934_ (.A_N(_2117_),
    .B(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__clkbuf_1 _3935_ (.A(_2123_),
    .X(_0557_));
 sky130_fd_sc_hd__xor2_1 _3936_ (.A(net136),
    .B(_2121_),
    .X(_0556_));
 sky130_fd_sc_hd__and3_1 _3937_ (.A(\output_c[15][16] ),
    .B(_2112_),
    .C(_2113_),
    .X(_2124_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(net382),
    .B(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__nor2_1 _3939_ (.A(_2121_),
    .B(_2125_),
    .Y(_0555_));
 sky130_fd_sc_hd__buf_1 _3940_ (.A(_2113_),
    .X(_2126_));
 sky130_fd_sc_hd__a21o_1 _3941_ (.A1(_2112_),
    .A2(_2126_),
    .B1(\output_c[15][16] ),
    .X(_2127_));
 sky130_fd_sc_hd__and2b_1 _3942_ (.A_N(_2124_),
    .B(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _3943_ (.A(_2128_),
    .X(_0554_));
 sky130_fd_sc_hd__and3_1 _3944_ (.A(\output_c[15][12] ),
    .B(_2096_),
    .C(_2097_),
    .X(_2129_));
 sky130_fd_sc_hd__and3_1 _3945_ (.A(\output_c[15][14] ),
    .B(\output_c[15][13] ),
    .C(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__xor2_1 _3946_ (.A(net64),
    .B(_2130_),
    .X(_0553_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3947_ (.A(_2126_),
    .X(_2131_));
 sky130_fd_sc_hd__a21oi_1 _3948_ (.A1(_2098_),
    .A2(_2131_),
    .B1(net344),
    .Y(_2132_));
 sky130_fd_sc_hd__nor2_1 _3949_ (.A(_2130_),
    .B(_2132_),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_1 _3950_ (.A(net311),
    .B(_2129_),
    .Y(_2133_));
 sky130_fd_sc_hd__a21oi_1 _3951_ (.A1(_2098_),
    .A2(_2131_),
    .B1(_2133_),
    .Y(_0551_));
 sky130_fd_sc_hd__and2_1 _3952_ (.A(_2097_),
    .B(_2126_),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_1 _3953_ (.A(net420),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__nor2_1 _3954_ (.A(_2129_),
    .B(_2135_),
    .Y(_0550_));
 sky130_fd_sc_hd__and3_1 _3955_ (.A(\output_c[15][9] ),
    .B(\output_c[15][8] ),
    .C(_2113_),
    .X(_2136_));
 sky130_fd_sc_hd__a21oi_1 _3956_ (.A1(\output_c[15][10] ),
    .A2(_2136_),
    .B1(net115),
    .Y(_2137_));
 sky130_fd_sc_hd__nor2_1 _3957_ (.A(_2134_),
    .B(net116),
    .Y(_0549_));
 sky130_fd_sc_hd__xor2_1 _3958_ (.A(net122),
    .B(_2136_),
    .X(_0548_));
 sky130_fd_sc_hd__a21oi_1 _3959_ (.A1(net272),
    .A2(_2131_),
    .B1(net405),
    .Y(_2138_));
 sky130_fd_sc_hd__nor2_1 _3960_ (.A(_2136_),
    .B(_2138_),
    .Y(_0547_));
 sky130_fd_sc_hd__xor2_1 _3961_ (.A(net272),
    .B(_2131_),
    .X(_0546_));
 sky130_fd_sc_hd__buf_1 _3962_ (.A(_2093_),
    .X(_2139_));
 sky130_fd_sc_hd__and3_1 _3963_ (.A(\output_c[15][5] ),
    .B(_2103_),
    .C(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__a21o_1 _3964_ (.A1(\output_c[15][6] ),
    .A2(_2140_),
    .B1(\output_c[15][7] ),
    .X(_2141_));
 sky130_fd_sc_hd__and2b_1 _3965_ (.A_N(_2126_),
    .B(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__clkbuf_1 _3966_ (.A(_2142_),
    .X(_0545_));
 sky130_fd_sc_hd__xor2_1 _3967_ (.A(net427),
    .B(_2140_),
    .X(_0544_));
 sky130_fd_sc_hd__a21oi_1 _3968_ (.A1(_2103_),
    .A2(_2139_),
    .B1(net470),
    .Y(_2143_));
 sky130_fd_sc_hd__nor2_1 _3969_ (.A(_2140_),
    .B(_2143_),
    .Y(_0543_));
 sky130_fd_sc_hd__xor2_1 _3970_ (.A(_2103_),
    .B(_2139_),
    .X(_0542_));
 sky130_fd_sc_hd__and3_1 _3971_ (.A(\output_c[15][1] ),
    .B(_1905_),
    .C(_2091_),
    .X(_2144_));
 sky130_fd_sc_hd__and2_1 _3972_ (.A(net421),
    .B(_2144_),
    .X(_2145_));
 sky130_fd_sc_hd__o21ba_1 _3973_ (.A1(net255),
    .A2(_2145_),
    .B1_N(_2139_),
    .X(_0541_));
 sky130_fd_sc_hd__nor2_1 _3974_ (.A(net421),
    .B(_2144_),
    .Y(_2146_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_2145_),
    .B(_2146_),
    .Y(_0540_));
 sky130_fd_sc_hd__a21oi_1 _3976_ (.A1(_1150_),
    .A2(_2091_),
    .B1(net320),
    .Y(_2147_));
 sky130_fd_sc_hd__nor2_1 _3977_ (.A(_2144_),
    .B(_2147_),
    .Y(_0539_));
 sky130_fd_sc_hd__and3_1 _3978_ (.A(_1348_),
    .B(\input_a[15] ),
    .C(_1911_),
    .X(_2148_));
 sky130_fd_sc_hd__o2bb2a_1 _3979_ (.A1_N(_1910_),
    .A2_N(_2091_),
    .B1(_2148_),
    .B2(net225),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(\input_a[14][0] ),
    .A1(_2048_),
    .S(_1220_),
    .X(_2149_));
 sky130_fd_sc_hd__clkbuf_1 _3981_ (.A(_2149_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_1 _3982_ (.A(_1345_),
    .X(_2150_));
 sky130_fd_sc_hd__and2_1 _3983_ (.A(\output_c[14][0] ),
    .B(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__buf_1 _3984_ (.A(_2151_),
    .X(net3));
 sky130_fd_sc_hd__and2_1 _3985_ (.A(\output_c[14][1] ),
    .B(_2150_),
    .X(_2152_));
 sky130_fd_sc_hd__buf_1 _3986_ (.A(_2152_),
    .X(net14));
 sky130_fd_sc_hd__and2_1 _3987_ (.A(_1076_),
    .B(_1150_),
    .X(_2153_));
 sky130_fd_sc_hd__buf_1 _3988_ (.A(_2153_),
    .X(net25));
 sky130_fd_sc_hd__and2_1 _3989_ (.A(\output_c[14][3] ),
    .B(_2150_),
    .X(_2154_));
 sky130_fd_sc_hd__buf_1 _3990_ (.A(_2154_),
    .X(net28));
 sky130_fd_sc_hd__buf_1 _3991_ (.A(_1143_),
    .X(_2155_));
 sky130_fd_sc_hd__buf_1 _3992_ (.A(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__and2_1 _3993_ (.A(_1135_),
    .B(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__buf_1 _3994_ (.A(_2157_),
    .X(net29));
 sky130_fd_sc_hd__and2_1 _3995_ (.A(_1134_),
    .B(_2156_),
    .X(_2158_));
 sky130_fd_sc_hd__buf_1 _3996_ (.A(_2158_),
    .X(net30));
 sky130_fd_sc_hd__and2_1 _3997_ (.A(\output_c[14][6] ),
    .B(_2156_),
    .X(_2159_));
 sky130_fd_sc_hd__buf_1 _3998_ (.A(_2159_),
    .X(net31));
 sky130_fd_sc_hd__and2_1 _3999_ (.A(\output_c[14][7] ),
    .B(_2156_),
    .X(_2160_));
 sky130_fd_sc_hd__buf_1 _4000_ (.A(_2160_),
    .X(net32));
 sky130_fd_sc_hd__buf_1 _4001_ (.A(_2155_),
    .X(_2161_));
 sky130_fd_sc_hd__and2_1 _4002_ (.A(\output_c[14][8] ),
    .B(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__buf_1 _4003_ (.A(_2162_),
    .X(net33));
 sky130_fd_sc_hd__and2_1 _4004_ (.A(_1128_),
    .B(_2161_),
    .X(_2163_));
 sky130_fd_sc_hd__buf_1 _4005_ (.A(_2163_),
    .X(net34));
 sky130_fd_sc_hd__and2_1 _4006_ (.A(\output_c[14][10] ),
    .B(_2161_),
    .X(_2164_));
 sky130_fd_sc_hd__buf_1 _4007_ (.A(_2164_),
    .X(net4));
 sky130_fd_sc_hd__and2_1 _4008_ (.A(\output_c[14][11] ),
    .B(_2161_),
    .X(_2165_));
 sky130_fd_sc_hd__buf_1 _4009_ (.A(_2165_),
    .X(net5));
 sky130_fd_sc_hd__buf_1 _4010_ (.A(_2155_),
    .X(_2166_));
 sky130_fd_sc_hd__and2_1 _4011_ (.A(\output_c[14][12] ),
    .B(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__buf_1 _4012_ (.A(_2167_),
    .X(net6));
 sky130_fd_sc_hd__and2_1 _4013_ (.A(_1122_),
    .B(_2166_),
    .X(_2168_));
 sky130_fd_sc_hd__buf_1 _4014_ (.A(_2168_),
    .X(net7));
 sky130_fd_sc_hd__and2_1 _4015_ (.A(\output_c[14][14] ),
    .B(_2166_),
    .X(_2169_));
 sky130_fd_sc_hd__clkbuf_1 _4016_ (.A(_2169_),
    .X(net8));
 sky130_fd_sc_hd__and2_1 _4017_ (.A(\output_c[14][15] ),
    .B(_2166_),
    .X(_2170_));
 sky130_fd_sc_hd__buf_1 _4018_ (.A(_2170_),
    .X(net9));
 sky130_fd_sc_hd__buf_1 _4019_ (.A(_2155_),
    .X(_2171_));
 sky130_fd_sc_hd__and2_1 _4020_ (.A(\output_c[14][16] ),
    .B(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__buf_1 _4021_ (.A(_2172_),
    .X(net10));
 sky130_fd_sc_hd__and2_1 _4022_ (.A(_1113_),
    .B(_2171_),
    .X(_2173_));
 sky130_fd_sc_hd__buf_1 _4023_ (.A(_2173_),
    .X(net11));
 sky130_fd_sc_hd__and2_1 _4024_ (.A(\output_c[14][18] ),
    .B(_2171_),
    .X(_2174_));
 sky130_fd_sc_hd__buf_1 _4025_ (.A(_2174_),
    .X(net12));
 sky130_fd_sc_hd__and2_1 _4026_ (.A(\output_c[14][19] ),
    .B(_2171_),
    .X(_2175_));
 sky130_fd_sc_hd__buf_1 _4027_ (.A(_2175_),
    .X(net13));
 sky130_fd_sc_hd__buf_1 _4028_ (.A(_1144_),
    .X(_2176_));
 sky130_fd_sc_hd__and2_1 _4029_ (.A(_1100_),
    .B(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__buf_1 _4030_ (.A(_2177_),
    .X(net15));
 sky130_fd_sc_hd__and2_1 _4031_ (.A(_1099_),
    .B(_2176_),
    .X(_2178_));
 sky130_fd_sc_hd__buf_1 _4032_ (.A(_2178_),
    .X(net16));
 sky130_fd_sc_hd__and2_1 _4033_ (.A(\output_c[14][22] ),
    .B(_2176_),
    .X(_2179_));
 sky130_fd_sc_hd__buf_1 _4034_ (.A(_2179_),
    .X(net17));
 sky130_fd_sc_hd__and2_1 _4035_ (.A(\output_c[14][23] ),
    .B(_2176_),
    .X(_2180_));
 sky130_fd_sc_hd__buf_1 _4036_ (.A(_2180_),
    .X(net18));
 sky130_fd_sc_hd__and2_1 _4037_ (.A(\output_c[14][24] ),
    .B(_2150_),
    .X(_2181_));
 sky130_fd_sc_hd__buf_1 _4038_ (.A(_2181_),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _4039_ (.A(_1144_),
    .X(_2182_));
 sky130_fd_sc_hd__and2_1 _4040_ (.A(_1091_),
    .B(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__buf_1 _4041_ (.A(_2183_),
    .X(net20));
 sky130_fd_sc_hd__and2_1 _4042_ (.A(\output_c[14][26] ),
    .B(_2182_),
    .X(_2184_));
 sky130_fd_sc_hd__buf_1 _4043_ (.A(_2184_),
    .X(net21));
 sky130_fd_sc_hd__and2_1 _4044_ (.A(\output_c[14][27] ),
    .B(_2182_),
    .X(_2185_));
 sky130_fd_sc_hd__buf_1 _4045_ (.A(_2185_),
    .X(net22));
 sky130_fd_sc_hd__and2_1 _4046_ (.A(\output_c[14][28] ),
    .B(_2182_),
    .X(_2186_));
 sky130_fd_sc_hd__buf_1 _4047_ (.A(_2186_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _4048_ (.A(\output_c[14][29] ),
    .B(_1156_),
    .X(_2187_));
 sky130_fd_sc_hd__buf_1 _4049_ (.A(_2187_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _4050_ (.A(\output_c[14][30] ),
    .B(_1156_),
    .X(_2188_));
 sky130_fd_sc_hd__buf_1 _4051_ (.A(_2188_),
    .X(net26));
 sky130_fd_sc_hd__and2_1 _4052_ (.A(\output_c[14][31] ),
    .B(_1156_),
    .X(_2189_));
 sky130_fd_sc_hd__buf_1 _4053_ (.A(_2189_),
    .X(net27));
 sky130_fd_sc_hd__nand2_1 _4054_ (.A(_2042_),
    .B(_2045_),
    .Y(_0001_));
 sky130_fd_sc_hd__xnor2_1 _4055_ (.A(_2055_),
    .B(_2079_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand3_1 _4056_ (.A(_2050_),
    .B(_2052_),
    .C(_2055_),
    .Y(_2190_));
 sky130_fd_sc_hd__a21o_1 _4057_ (.A1(_2056_),
    .A2(_2190_),
    .B1(_2069_),
    .X(_0003_));
 sky130_fd_sc_hd__clkbuf_2 _4058_ (.A(net2),
    .X(_2191_));
 sky130_fd_sc_hd__buf_1 _4059_ (.A(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4060_ (.A(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_2 _4061_ (.A(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__inv_2 _4062_ (.A(_2194_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _4063_ (.A(_2194_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _4064_ (.A(_2194_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _4065_ (.A(_2194_),
    .Y(_0007_));
 sky130_fd_sc_hd__clkbuf_2 _4066_ (.A(_2193_),
    .X(_2195_));
 sky130_fd_sc_hd__inv_2 _4067_ (.A(_2195_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _4068_ (.A(_2195_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _4069_ (.A(_2195_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _4070_ (.A(_2195_),
    .Y(_0011_));
 sky130_fd_sc_hd__clkbuf_2 _4071_ (.A(_2193_),
    .X(_2196_));
 sky130_fd_sc_hd__inv_2 _4072_ (.A(_2196_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _4073_ (.A(_2196_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _4074_ (.A(_2196_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _4075_ (.A(_2196_),
    .Y(_0015_));
 sky130_fd_sc_hd__buf_1 _4076_ (.A(_2191_),
    .X(_2197_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4077_ (.A(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__clkbuf_2 _4078_ (.A(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__inv_2 _4079_ (.A(_2199_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _4080_ (.A(_2199_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _4081_ (.A(_2199_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _4082_ (.A(_2199_),
    .Y(_0019_));
 sky130_fd_sc_hd__clkbuf_2 _4083_ (.A(_2198_),
    .X(_2200_));
 sky130_fd_sc_hd__inv_2 _4084_ (.A(_2200_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _4085_ (.A(_2200_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _4086_ (.A(_2200_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _4087_ (.A(_2200_),
    .Y(_0023_));
 sky130_fd_sc_hd__clkbuf_2 _4088_ (.A(_2198_),
    .X(_2201_));
 sky130_fd_sc_hd__inv_2 _4089_ (.A(_2201_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _4090_ (.A(_2201_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _4091_ (.A(_2201_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _4092_ (.A(_2201_),
    .Y(_0027_));
 sky130_fd_sc_hd__clkbuf_2 _4093_ (.A(_2198_),
    .X(_2202_));
 sky130_fd_sc_hd__inv_2 _4094_ (.A(_2202_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _4095_ (.A(_2202_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _4096_ (.A(_2202_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _4097_ (.A(_2202_),
    .Y(_0031_));
 sky130_fd_sc_hd__clkbuf_2 _4098_ (.A(_2197_),
    .X(_2203_));
 sky130_fd_sc_hd__clkbuf_2 _4099_ (.A(_2203_),
    .X(_2204_));
 sky130_fd_sc_hd__inv_2 _4100_ (.A(_2204_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _4101_ (.A(_2204_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _4102_ (.A(_2204_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _4103_ (.A(_2204_),
    .Y(_0035_));
 sky130_fd_sc_hd__clkbuf_2 _4104_ (.A(_2203_),
    .X(_2205_));
 sky130_fd_sc_hd__inv_2 _4105_ (.A(_2205_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _4106_ (.A(_2205_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _4107_ (.A(_2205_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _4108_ (.A(_2205_),
    .Y(_0039_));
 sky130_fd_sc_hd__clkbuf_2 _4109_ (.A(_2203_),
    .X(_2206_));
 sky130_fd_sc_hd__inv_2 _4110_ (.A(_2206_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _4111_ (.A(_2206_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _4112_ (.A(_2206_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _4113_ (.A(_2206_),
    .Y(_0043_));
 sky130_fd_sc_hd__clkbuf_2 _4114_ (.A(_2203_),
    .X(_2207_));
 sky130_fd_sc_hd__inv_2 _4115_ (.A(_2207_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _4116_ (.A(_2207_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _4117_ (.A(_2207_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _4118_ (.A(_2207_),
    .Y(_0047_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4119_ (.A(_2192_),
    .X(_2208_));
 sky130_fd_sc_hd__buf_1 _4120_ (.A(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__clkbuf_2 _4121_ (.A(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__inv_2 _4122_ (.A(_2210_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _4123_ (.A(_2210_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _4124_ (.A(_2210_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _4125_ (.A(_2210_),
    .Y(_0051_));
 sky130_fd_sc_hd__clkbuf_2 _4126_ (.A(_2209_),
    .X(_2211_));
 sky130_fd_sc_hd__inv_2 _4127_ (.A(_2211_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _4128_ (.A(_2211_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _4129_ (.A(_2211_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _4130_ (.A(_2211_),
    .Y(_0055_));
 sky130_fd_sc_hd__clkbuf_2 _4131_ (.A(_2209_),
    .X(_2212_));
 sky130_fd_sc_hd__inv_2 _4132_ (.A(_2212_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _4133_ (.A(_2212_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _4134_ (.A(_2212_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _4135_ (.A(_2212_),
    .Y(_0059_));
 sky130_fd_sc_hd__clkbuf_2 _4136_ (.A(_2209_),
    .X(_2213_));
 sky130_fd_sc_hd__inv_2 _4137_ (.A(_2213_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _4138_ (.A(_2213_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _4139_ (.A(_2213_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _4140_ (.A(_2213_),
    .Y(_0063_));
 sky130_fd_sc_hd__buf_1 _4141_ (.A(_2208_),
    .X(_2214_));
 sky130_fd_sc_hd__clkbuf_2 _4142_ (.A(_2214_),
    .X(_2215_));
 sky130_fd_sc_hd__inv_2 _4143_ (.A(_2215_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _4144_ (.A(_2215_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _4145_ (.A(_2215_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _4146_ (.A(_2215_),
    .Y(_0067_));
 sky130_fd_sc_hd__clkbuf_2 _4147_ (.A(_2214_),
    .X(_2216_));
 sky130_fd_sc_hd__inv_2 _4148_ (.A(_2216_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _4149_ (.A(_2216_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _4150_ (.A(_2216_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _4151_ (.A(_2216_),
    .Y(_0071_));
 sky130_fd_sc_hd__clkbuf_2 _4152_ (.A(_2214_),
    .X(_2217_));
 sky130_fd_sc_hd__inv_2 _4153_ (.A(_2217_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _4154_ (.A(_2217_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _4155_ (.A(_2217_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _4156_ (.A(_2217_),
    .Y(_0075_));
 sky130_fd_sc_hd__clkbuf_2 _4157_ (.A(_2214_),
    .X(_2218_));
 sky130_fd_sc_hd__inv_2 _4158_ (.A(_2218_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _4159_ (.A(_2218_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _4160_ (.A(_2218_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _4161_ (.A(_2218_),
    .Y(_0079_));
 sky130_fd_sc_hd__buf_1 _4162_ (.A(_2208_),
    .X(_2219_));
 sky130_fd_sc_hd__clkbuf_2 _4163_ (.A(_2219_),
    .X(_2220_));
 sky130_fd_sc_hd__inv_2 _4164_ (.A(_2220_),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _4165_ (.A(_2220_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _4166_ (.A(_2220_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _4167_ (.A(_2220_),
    .Y(_0083_));
 sky130_fd_sc_hd__clkbuf_2 _4168_ (.A(_2219_),
    .X(_2221_));
 sky130_fd_sc_hd__inv_2 _4169_ (.A(_2221_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _4170_ (.A(_2221_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _4171_ (.A(_2221_),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _4172_ (.A(_2221_),
    .Y(_0087_));
 sky130_fd_sc_hd__clkbuf_2 _4173_ (.A(_2219_),
    .X(_2222_));
 sky130_fd_sc_hd__inv_2 _4174_ (.A(_2222_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _4175_ (.A(_2222_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _4176_ (.A(_2222_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _4177_ (.A(_2222_),
    .Y(_0091_));
 sky130_fd_sc_hd__clkbuf_2 _4178_ (.A(_2219_),
    .X(_2223_));
 sky130_fd_sc_hd__inv_2 _4179_ (.A(_2223_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _4180_ (.A(_2223_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _4181_ (.A(_2223_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _4182_ (.A(_2223_),
    .Y(_0095_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4183_ (.A(_2208_),
    .X(_2224_));
 sky130_fd_sc_hd__clkbuf_2 _4184_ (.A(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(_2225_),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _4186_ (.A(_2225_),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _4187_ (.A(_2225_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _4188_ (.A(_2225_),
    .Y(_0099_));
 sky130_fd_sc_hd__clkbuf_2 _4189_ (.A(_2224_),
    .X(_2226_));
 sky130_fd_sc_hd__inv_2 _4190_ (.A(_2226_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _4191_ (.A(_2226_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _4192_ (.A(_2226_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _4193_ (.A(_2226_),
    .Y(_0103_));
 sky130_fd_sc_hd__clkbuf_2 _4194_ (.A(_2224_),
    .X(_2227_));
 sky130_fd_sc_hd__inv_2 _4195_ (.A(_2227_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _4196_ (.A(_2227_),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(_2227_),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _4198_ (.A(_2227_),
    .Y(_0107_));
 sky130_fd_sc_hd__clkbuf_2 _4199_ (.A(_2224_),
    .X(_2228_));
 sky130_fd_sc_hd__inv_2 _4200_ (.A(_2228_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _4201_ (.A(_2228_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _4202_ (.A(_2228_),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _4203_ (.A(_2228_),
    .Y(_0111_));
 sky130_fd_sc_hd__clkbuf_2 _4204_ (.A(net2),
    .X(_2229_));
 sky130_fd_sc_hd__buf_1 _4205_ (.A(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__buf_1 _4206_ (.A(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__clkbuf_2 _4207_ (.A(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__inv_2 _4208_ (.A(_2232_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _4209_ (.A(_2232_),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _4210_ (.A(_2232_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _4211_ (.A(_2232_),
    .Y(_0115_));
 sky130_fd_sc_hd__clkbuf_2 _4212_ (.A(_2231_),
    .X(_2233_));
 sky130_fd_sc_hd__inv_2 _4213_ (.A(_2233_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _4214_ (.A(_2233_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _4215_ (.A(_2233_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _4216_ (.A(_2233_),
    .Y(_0119_));
 sky130_fd_sc_hd__clkbuf_2 _4217_ (.A(_2231_),
    .X(_2234_));
 sky130_fd_sc_hd__inv_2 _4218_ (.A(_2234_),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _4219_ (.A(_2234_),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _4220_ (.A(_2234_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _4221_ (.A(_2234_),
    .Y(_0123_));
 sky130_fd_sc_hd__clkbuf_2 _4222_ (.A(_2231_),
    .X(_2235_));
 sky130_fd_sc_hd__inv_2 _4223_ (.A(_2235_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _4224_ (.A(_2235_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _4225_ (.A(_2235_),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _4226_ (.A(_2235_),
    .Y(_0127_));
 sky130_fd_sc_hd__buf_1 _4227_ (.A(_2230_),
    .X(_2236_));
 sky130_fd_sc_hd__clkbuf_2 _4228_ (.A(_2236_),
    .X(_2237_));
 sky130_fd_sc_hd__inv_2 _4229_ (.A(_2237_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _4230_ (.A(_2237_),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _4231_ (.A(_2237_),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _4232_ (.A(_2237_),
    .Y(_0131_));
 sky130_fd_sc_hd__clkbuf_2 _4233_ (.A(_2236_),
    .X(_2238_));
 sky130_fd_sc_hd__inv_2 _4234_ (.A(_2238_),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _4235_ (.A(_2238_),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _4236_ (.A(_2238_),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _4237_ (.A(_2238_),
    .Y(_0135_));
 sky130_fd_sc_hd__clkbuf_2 _4238_ (.A(_2236_),
    .X(_2239_));
 sky130_fd_sc_hd__inv_2 _4239_ (.A(_2239_),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _4240_ (.A(_2239_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _4241_ (.A(_2239_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _4242_ (.A(_2239_),
    .Y(_0139_));
 sky130_fd_sc_hd__clkbuf_2 _4243_ (.A(_2236_),
    .X(_2240_));
 sky130_fd_sc_hd__inv_2 _4244_ (.A(_2240_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _4245_ (.A(_2240_),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _4246_ (.A(_2240_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _4247_ (.A(_2240_),
    .Y(_0143_));
 sky130_fd_sc_hd__buf_1 _4248_ (.A(_2230_),
    .X(_2241_));
 sky130_fd_sc_hd__clkbuf_2 _4249_ (.A(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__inv_2 _4250_ (.A(_2242_),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _4251_ (.A(_2242_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _4252_ (.A(_2242_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _4253_ (.A(_2242_),
    .Y(_0147_));
 sky130_fd_sc_hd__clkbuf_2 _4254_ (.A(_2241_),
    .X(_2243_));
 sky130_fd_sc_hd__inv_2 _4255_ (.A(_2243_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _4256_ (.A(_2243_),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _4257_ (.A(_2243_),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _4258_ (.A(_2243_),
    .Y(_0151_));
 sky130_fd_sc_hd__clkbuf_2 _4259_ (.A(_2241_),
    .X(_2244_));
 sky130_fd_sc_hd__inv_2 _4260_ (.A(_2244_),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _4261_ (.A(_2244_),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _4262_ (.A(_2244_),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _4263_ (.A(_2244_),
    .Y(_0155_));
 sky130_fd_sc_hd__clkbuf_2 _4264_ (.A(_2241_),
    .X(_2245_));
 sky130_fd_sc_hd__inv_2 _4265_ (.A(_2245_),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _4266_ (.A(_2245_),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _4267_ (.A(_2245_),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _4268_ (.A(_2245_),
    .Y(_0159_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4269_ (.A(_2230_),
    .X(_2246_));
 sky130_fd_sc_hd__clkbuf_2 _4270_ (.A(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__inv_2 _4271_ (.A(_2247_),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _4272_ (.A(_2247_),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _4273_ (.A(_2247_),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _4274_ (.A(_2247_),
    .Y(_0163_));
 sky130_fd_sc_hd__clkbuf_2 _4275_ (.A(_2246_),
    .X(_2248_));
 sky130_fd_sc_hd__inv_2 _4276_ (.A(_2248_),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _4277_ (.A(_2248_),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _4278_ (.A(_2248_),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _4279_ (.A(_2248_),
    .Y(_0167_));
 sky130_fd_sc_hd__clkbuf_2 _4280_ (.A(_2246_),
    .X(_2249_));
 sky130_fd_sc_hd__inv_2 _4281_ (.A(_2249_),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _4282_ (.A(_2249_),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _4283_ (.A(_2249_),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _4284_ (.A(_2249_),
    .Y(_0171_));
 sky130_fd_sc_hd__clkbuf_2 _4285_ (.A(_2246_),
    .X(_2250_));
 sky130_fd_sc_hd__inv_2 _4286_ (.A(_2250_),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _4287_ (.A(_2250_),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _4288_ (.A(_2250_),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _4289_ (.A(_2250_),
    .Y(_0175_));
 sky130_fd_sc_hd__buf_1 _4290_ (.A(_2229_),
    .X(_2251_));
 sky130_fd_sc_hd__buf_1 _4291_ (.A(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__clkbuf_2 _4292_ (.A(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__inv_2 _4293_ (.A(_2253_),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _4294_ (.A(_2253_),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _4295_ (.A(_2253_),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _4296_ (.A(_2253_),
    .Y(_0179_));
 sky130_fd_sc_hd__clkbuf_2 _4297_ (.A(_2252_),
    .X(_2254_));
 sky130_fd_sc_hd__inv_2 _4298_ (.A(_2254_),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _4299_ (.A(_2254_),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _4300_ (.A(_2254_),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _4301_ (.A(_2254_),
    .Y(_0183_));
 sky130_fd_sc_hd__buf_2 _4302_ (.A(_2252_),
    .X(_2255_));
 sky130_fd_sc_hd__inv_2 _4303_ (.A(_2255_),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _4304_ (.A(_2255_),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _4305_ (.A(_2255_),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _4306_ (.A(_2255_),
    .Y(_0187_));
 sky130_fd_sc_hd__clkbuf_2 _4307_ (.A(_2252_),
    .X(_2256_));
 sky130_fd_sc_hd__inv_2 _4308_ (.A(_2256_),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _4309_ (.A(_2256_),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _4310_ (.A(_2256_),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _4311_ (.A(_2256_),
    .Y(_0191_));
 sky130_fd_sc_hd__buf_1 _4312_ (.A(_2251_),
    .X(_2257_));
 sky130_fd_sc_hd__clkbuf_2 _4313_ (.A(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__inv_2 _4314_ (.A(_2258_),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _4315_ (.A(_2258_),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _4316_ (.A(_2258_),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _4317_ (.A(_2258_),
    .Y(_0195_));
 sky130_fd_sc_hd__clkbuf_2 _4318_ (.A(_2257_),
    .X(_2259_));
 sky130_fd_sc_hd__inv_2 _4319_ (.A(_2259_),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _4320_ (.A(_2259_),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _4321_ (.A(_2259_),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _4322_ (.A(_2259_),
    .Y(_0199_));
 sky130_fd_sc_hd__clkbuf_2 _4323_ (.A(_2257_),
    .X(_2260_));
 sky130_fd_sc_hd__inv_2 _4324_ (.A(_2260_),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _4325_ (.A(_2260_),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _4326_ (.A(_2260_),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _4327_ (.A(_2260_),
    .Y(_0203_));
 sky130_fd_sc_hd__clkbuf_2 _4328_ (.A(_2257_),
    .X(_2261_));
 sky130_fd_sc_hd__inv_2 _4329_ (.A(_2261_),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _4330_ (.A(_2261_),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _4331_ (.A(_2261_),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _4332_ (.A(_2261_),
    .Y(_0207_));
 sky130_fd_sc_hd__buf_1 _4333_ (.A(_2251_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_2 _4334_ (.A(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__inv_2 _4335_ (.A(_2263_),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _4336_ (.A(_2263_),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _4337_ (.A(_2263_),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _4338_ (.A(_2263_),
    .Y(_0211_));
 sky130_fd_sc_hd__clkbuf_2 _4339_ (.A(_2262_),
    .X(_2264_));
 sky130_fd_sc_hd__inv_2 _4340_ (.A(_2264_),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _4341_ (.A(_2264_),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _4342_ (.A(_2264_),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _4343_ (.A(_2264_),
    .Y(_0215_));
 sky130_fd_sc_hd__clkbuf_2 _4344_ (.A(_2262_),
    .X(_2265_));
 sky130_fd_sc_hd__inv_2 _4345_ (.A(_2265_),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _4346_ (.A(_2265_),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_2 _4347_ (.A(_2265_),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _4348_ (.A(_2265_),
    .Y(_0219_));
 sky130_fd_sc_hd__clkbuf_2 _4349_ (.A(_2262_),
    .X(_2266_));
 sky130_fd_sc_hd__inv_2 _4350_ (.A(_2266_),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _4351_ (.A(_2266_),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _4352_ (.A(_2266_),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _4353_ (.A(_2266_),
    .Y(_0223_));
 sky130_fd_sc_hd__buf_1 _4354_ (.A(_2251_),
    .X(_2267_));
 sky130_fd_sc_hd__clkbuf_2 _4355_ (.A(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__inv_2 _4356_ (.A(_2268_),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _4357_ (.A(_2268_),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _4358_ (.A(_2268_),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _4359_ (.A(_2268_),
    .Y(_0227_));
 sky130_fd_sc_hd__clkbuf_2 _4360_ (.A(_2267_),
    .X(_2269_));
 sky130_fd_sc_hd__inv_2 _4361_ (.A(_2269_),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _4362_ (.A(_2269_),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_2 _4363_ (.A(_2269_),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_2 _4364_ (.A(_2269_),
    .Y(_0231_));
 sky130_fd_sc_hd__clkbuf_2 _4365_ (.A(_2267_),
    .X(_2270_));
 sky130_fd_sc_hd__inv_2 _4366_ (.A(_2270_),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _4367_ (.A(_2270_),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _4368_ (.A(_2270_),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _4369_ (.A(_2270_),
    .Y(_0235_));
 sky130_fd_sc_hd__clkbuf_2 _4370_ (.A(_2267_),
    .X(_2271_));
 sky130_fd_sc_hd__inv_2 _4371_ (.A(_2271_),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _4372_ (.A(_2271_),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _4373_ (.A(_2271_),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _4374_ (.A(_2271_),
    .Y(_0239_));
 sky130_fd_sc_hd__clkbuf_2 _4375_ (.A(_2229_),
    .X(_2272_));
 sky130_fd_sc_hd__buf_1 _4376_ (.A(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__clkbuf_2 _4377_ (.A(_2273_),
    .X(_2274_));
 sky130_fd_sc_hd__inv_2 _4378_ (.A(_2274_),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _4379_ (.A(_2274_),
    .Y(_0241_));
 sky130_fd_sc_hd__inv_2 _4380_ (.A(_2274_),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _4381_ (.A(_2274_),
    .Y(_0243_));
 sky130_fd_sc_hd__clkbuf_2 _4382_ (.A(_2273_),
    .X(_2275_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(_2275_),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _4384_ (.A(_2275_),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _4385_ (.A(_2275_),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _4386_ (.A(_2275_),
    .Y(_0247_));
 sky130_fd_sc_hd__clkbuf_2 _4387_ (.A(_2273_),
    .X(_2276_));
 sky130_fd_sc_hd__inv_2 _4388_ (.A(_2276_),
    .Y(_0248_));
 sky130_fd_sc_hd__inv_2 _4389_ (.A(_2276_),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_2 _4390_ (.A(_2276_),
    .Y(_0250_));
 sky130_fd_sc_hd__inv_2 _4391_ (.A(_2276_),
    .Y(_0251_));
 sky130_fd_sc_hd__clkbuf_2 _4392_ (.A(_2273_),
    .X(_2277_));
 sky130_fd_sc_hd__inv_2 _4393_ (.A(_2277_),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _4394_ (.A(_2277_),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _4395_ (.A(_2277_),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _4396_ (.A(_2277_),
    .Y(_0255_));
 sky130_fd_sc_hd__buf_1 _4397_ (.A(_2272_),
    .X(_2278_));
 sky130_fd_sc_hd__clkbuf_2 _4398_ (.A(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__inv_2 _4399_ (.A(_2279_),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _4400_ (.A(_2279_),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_2 _4401_ (.A(_2279_),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_2 _4402_ (.A(_2279_),
    .Y(_0259_));
 sky130_fd_sc_hd__clkbuf_2 _4403_ (.A(_2278_),
    .X(_2280_));
 sky130_fd_sc_hd__inv_2 _4404_ (.A(_2280_),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _4405_ (.A(_2280_),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _4406_ (.A(_2280_),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _4407_ (.A(_2280_),
    .Y(_0263_));
 sky130_fd_sc_hd__clkbuf_2 _4408_ (.A(_2278_),
    .X(_2281_));
 sky130_fd_sc_hd__inv_2 _4409_ (.A(_2281_),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _4410_ (.A(_2281_),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_2 _4411_ (.A(_2281_),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _4412_ (.A(_2281_),
    .Y(_0267_));
 sky130_fd_sc_hd__clkbuf_2 _4413_ (.A(_2278_),
    .X(_2282_));
 sky130_fd_sc_hd__inv_2 _4414_ (.A(_2282_),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _4415_ (.A(_2282_),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _4416_ (.A(_2282_),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _4417_ (.A(_2282_),
    .Y(_0271_));
 sky130_fd_sc_hd__buf_1 _4418_ (.A(_2272_),
    .X(_2283_));
 sky130_fd_sc_hd__clkbuf_2 _4419_ (.A(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__inv_2 _4420_ (.A(_2284_),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _4421_ (.A(_2284_),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _4422_ (.A(_2284_),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _4423_ (.A(_2284_),
    .Y(_0275_));
 sky130_fd_sc_hd__clkbuf_2 _4424_ (.A(_2283_),
    .X(_2285_));
 sky130_fd_sc_hd__inv_2 _4425_ (.A(_2285_),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _4426_ (.A(_2285_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _4427_ (.A(_2285_),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _4428_ (.A(_2285_),
    .Y(_0279_));
 sky130_fd_sc_hd__buf_2 _4429_ (.A(_2283_),
    .X(_2286_));
 sky130_fd_sc_hd__inv_2 _4430_ (.A(_2286_),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _4431_ (.A(_2286_),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _4432_ (.A(_2286_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _4433_ (.A(_2286_),
    .Y(_0283_));
 sky130_fd_sc_hd__clkbuf_2 _4434_ (.A(_2283_),
    .X(_2287_));
 sky130_fd_sc_hd__inv_2 _4435_ (.A(_2287_),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _4436_ (.A(_2287_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _4437_ (.A(_2287_),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _4438_ (.A(_2287_),
    .Y(_0287_));
 sky130_fd_sc_hd__buf_1 _4439_ (.A(_2272_),
    .X(_2288_));
 sky130_fd_sc_hd__clkbuf_2 _4440_ (.A(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__inv_2 _4441_ (.A(_2289_),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _4442_ (.A(_2289_),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_2 _4443_ (.A(_2289_),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_2 _4444_ (.A(_2289_),
    .Y(_0291_));
 sky130_fd_sc_hd__clkbuf_2 _4445_ (.A(_2288_),
    .X(_2290_));
 sky130_fd_sc_hd__inv_2 _4446_ (.A(_2290_),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _4447_ (.A(_2290_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _4448_ (.A(_2290_),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_2 _4449_ (.A(_2290_),
    .Y(_0295_));
 sky130_fd_sc_hd__clkbuf_2 _4450_ (.A(_2288_),
    .X(_2291_));
 sky130_fd_sc_hd__inv_2 _4451_ (.A(_2291_),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_2 _4452_ (.A(_2291_),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _4453_ (.A(_2291_),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _4454_ (.A(_2291_),
    .Y(_0299_));
 sky130_fd_sc_hd__clkbuf_2 _4455_ (.A(_2288_),
    .X(_2292_));
 sky130_fd_sc_hd__inv_2 _4456_ (.A(_2292_),
    .Y(_0300_));
 sky130_fd_sc_hd__inv_2 _4457_ (.A(_2292_),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_2 _4458_ (.A(_2292_),
    .Y(_0302_));
 sky130_fd_sc_hd__inv_2 _4459_ (.A(_2292_),
    .Y(_0303_));
 sky130_fd_sc_hd__clkbuf_2 _4460_ (.A(_2229_),
    .X(_2293_));
 sky130_fd_sc_hd__clkbuf_2 _4461_ (.A(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__clkbuf_2 _4462_ (.A(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__inv_2 _4463_ (.A(_2295_),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _4464_ (.A(_2295_),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _4465_ (.A(_2295_),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _4466_ (.A(_2295_),
    .Y(_0307_));
 sky130_fd_sc_hd__clkbuf_2 _4467_ (.A(_2294_),
    .X(_2296_));
 sky130_fd_sc_hd__inv_2 _4468_ (.A(_2296_),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _4469_ (.A(_2296_),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _4470_ (.A(_2296_),
    .Y(_0310_));
 sky130_fd_sc_hd__inv_2 _4471_ (.A(_2296_),
    .Y(_0311_));
 sky130_fd_sc_hd__clkbuf_2 _4472_ (.A(_2294_),
    .X(_2297_));
 sky130_fd_sc_hd__inv_2 _4473_ (.A(_2297_),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _4474_ (.A(_2297_),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_2 _4475_ (.A(_2297_),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _4476_ (.A(_2297_),
    .Y(_0315_));
 sky130_fd_sc_hd__clkbuf_2 _4477_ (.A(_2294_),
    .X(_2298_));
 sky130_fd_sc_hd__inv_2 _4478_ (.A(_2298_),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _4479_ (.A(_2298_),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _4480_ (.A(_2298_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _4481_ (.A(_2298_),
    .Y(_0319_));
 sky130_fd_sc_hd__buf_1 _4482_ (.A(_2293_),
    .X(_2299_));
 sky130_fd_sc_hd__clkbuf_2 _4483_ (.A(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__inv_2 _4484_ (.A(_2300_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _4485_ (.A(_2300_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _4486_ (.A(_2300_),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _4487_ (.A(_2300_),
    .Y(_0323_));
 sky130_fd_sc_hd__clkbuf_2 _4488_ (.A(_2299_),
    .X(_2301_));
 sky130_fd_sc_hd__inv_2 _4489_ (.A(_2301_),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _4490_ (.A(_2301_),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _4491_ (.A(_2301_),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _4492_ (.A(_2301_),
    .Y(_0327_));
 sky130_fd_sc_hd__clkbuf_2 _4493_ (.A(_2299_),
    .X(_2302_));
 sky130_fd_sc_hd__inv_2 _4494_ (.A(_2302_),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _4495_ (.A(_2302_),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _4496_ (.A(_2302_),
    .Y(_0330_));
 sky130_fd_sc_hd__inv_2 _4497_ (.A(_2302_),
    .Y(_0331_));
 sky130_fd_sc_hd__clkbuf_2 _4498_ (.A(_2299_),
    .X(_2303_));
 sky130_fd_sc_hd__inv_2 _4499_ (.A(_2303_),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _4500_ (.A(_2303_),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _4501_ (.A(_2303_),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _4502_ (.A(_2303_),
    .Y(_0335_));
 sky130_fd_sc_hd__buf_1 _4503_ (.A(_2293_),
    .X(_2304_));
 sky130_fd_sc_hd__clkbuf_2 _4504_ (.A(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__inv_2 _4505_ (.A(_2305_),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _4506_ (.A(_2305_),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _4507_ (.A(_2305_),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _4508_ (.A(_2305_),
    .Y(_0339_));
 sky130_fd_sc_hd__clkbuf_2 _4509_ (.A(_2304_),
    .X(_2306_));
 sky130_fd_sc_hd__inv_2 _4510_ (.A(_2306_),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _4511_ (.A(_2306_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _4512_ (.A(_2306_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _4513_ (.A(_2306_),
    .Y(_0343_));
 sky130_fd_sc_hd__clkbuf_2 _4514_ (.A(_2304_),
    .X(_2307_));
 sky130_fd_sc_hd__inv_2 _4515_ (.A(_2307_),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _4516_ (.A(_2307_),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _4517_ (.A(_2307_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _4518_ (.A(_2307_),
    .Y(_0347_));
 sky130_fd_sc_hd__clkbuf_2 _4519_ (.A(_2304_),
    .X(_2308_));
 sky130_fd_sc_hd__inv_2 _4520_ (.A(_2308_),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _4521_ (.A(_2308_),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _4522_ (.A(_2308_),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_2 _4523_ (.A(_2308_),
    .Y(_0351_));
 sky130_fd_sc_hd__buf_1 _4524_ (.A(_2293_),
    .X(_2309_));
 sky130_fd_sc_hd__clkbuf_2 _4525_ (.A(_2309_),
    .X(_2310_));
 sky130_fd_sc_hd__inv_2 _4526_ (.A(_2310_),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _4527_ (.A(_2310_),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _4528_ (.A(_2310_),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _4529_ (.A(_2310_),
    .Y(_0355_));
 sky130_fd_sc_hd__clkbuf_2 _4530_ (.A(_2309_),
    .X(_2311_));
 sky130_fd_sc_hd__inv_2 _4531_ (.A(_2311_),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _4532_ (.A(_2311_),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _4533_ (.A(_2311_),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_2 _4534_ (.A(_2311_),
    .Y(_0359_));
 sky130_fd_sc_hd__clkbuf_2 _4535_ (.A(_2309_),
    .X(_2312_));
 sky130_fd_sc_hd__inv_2 _4536_ (.A(_2312_),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_2 _4537_ (.A(_2312_),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _4538_ (.A(_2312_),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _4539_ (.A(_2312_),
    .Y(_0363_));
 sky130_fd_sc_hd__clkbuf_2 _4540_ (.A(_2309_),
    .X(_2313_));
 sky130_fd_sc_hd__inv_2 _4541_ (.A(_2313_),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_2 _4542_ (.A(_2313_),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_2 _4543_ (.A(_2313_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _4544_ (.A(_2313_),
    .Y(_0367_));
 sky130_fd_sc_hd__clkbuf_2 _4545_ (.A(_2191_),
    .X(_2314_));
 sky130_fd_sc_hd__buf_1 _4546_ (.A(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__clkbuf_2 _4547_ (.A(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__inv_2 _4548_ (.A(_2316_),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _4549_ (.A(_2316_),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_2 _4550_ (.A(_2316_),
    .Y(_0370_));
 sky130_fd_sc_hd__inv_2 _4551_ (.A(_2316_),
    .Y(_0371_));
 sky130_fd_sc_hd__clkbuf_2 _4552_ (.A(_2315_),
    .X(_2317_));
 sky130_fd_sc_hd__inv_2 _4553_ (.A(_2317_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _4554_ (.A(_2317_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _4555_ (.A(_2317_),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _4556_ (.A(_2317_),
    .Y(_0375_));
 sky130_fd_sc_hd__clkbuf_2 _4557_ (.A(_2315_),
    .X(_2318_));
 sky130_fd_sc_hd__inv_2 _4558_ (.A(_2318_),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _4559_ (.A(_2318_),
    .Y(_0377_));
 sky130_fd_sc_hd__inv_2 _4560_ (.A(_2318_),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_2 _4561_ (.A(_2318_),
    .Y(_0379_));
 sky130_fd_sc_hd__clkbuf_2 _4562_ (.A(_2315_),
    .X(_2319_));
 sky130_fd_sc_hd__inv_2 _4563_ (.A(_2319_),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _4564_ (.A(_2319_),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_2 _4565_ (.A(_2319_),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_2 _4566_ (.A(_2319_),
    .Y(_0383_));
 sky130_fd_sc_hd__buf_1 _4567_ (.A(_2314_),
    .X(_2320_));
 sky130_fd_sc_hd__clkbuf_2 _4568_ (.A(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__inv_2 _4569_ (.A(_2321_),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_2 _4570_ (.A(_2321_),
    .Y(_0385_));
 sky130_fd_sc_hd__inv_2 _4571_ (.A(_2321_),
    .Y(_0386_));
 sky130_fd_sc_hd__inv_2 _4572_ (.A(_2321_),
    .Y(_0387_));
 sky130_fd_sc_hd__clkbuf_2 _4573_ (.A(_2320_),
    .X(_2322_));
 sky130_fd_sc_hd__inv_2 _4574_ (.A(_2322_),
    .Y(_0388_));
 sky130_fd_sc_hd__inv_2 _4575_ (.A(_2322_),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_2 _4576_ (.A(_2322_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _4577_ (.A(_2322_),
    .Y(_0391_));
 sky130_fd_sc_hd__clkbuf_2 _4578_ (.A(_2320_),
    .X(_2323_));
 sky130_fd_sc_hd__inv_2 _4579_ (.A(_2323_),
    .Y(_0392_));
 sky130_fd_sc_hd__inv_2 _4580_ (.A(_2323_),
    .Y(_0393_));
 sky130_fd_sc_hd__inv_2 _4581_ (.A(_2323_),
    .Y(_0394_));
 sky130_fd_sc_hd__inv_2 _4582_ (.A(_2323_),
    .Y(_0395_));
 sky130_fd_sc_hd__clkbuf_2 _4583_ (.A(_2320_),
    .X(_2324_));
 sky130_fd_sc_hd__inv_2 _4584_ (.A(_2324_),
    .Y(_0396_));
 sky130_fd_sc_hd__inv_2 _4585_ (.A(_2324_),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_2 _4586_ (.A(_2324_),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _4587_ (.A(_2324_),
    .Y(_0399_));
 sky130_fd_sc_hd__buf_1 _4588_ (.A(_2314_),
    .X(_2325_));
 sky130_fd_sc_hd__clkbuf_2 _4589_ (.A(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__inv_2 _4590_ (.A(_2326_),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_2 _4591_ (.A(_2326_),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _4592_ (.A(_2326_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _4593_ (.A(_2326_),
    .Y(_0403_));
 sky130_fd_sc_hd__clkbuf_2 _4594_ (.A(_2325_),
    .X(_2327_));
 sky130_fd_sc_hd__inv_2 _4595_ (.A(_2327_),
    .Y(_0404_));
 sky130_fd_sc_hd__inv_2 _4596_ (.A(_2327_),
    .Y(_0405_));
 sky130_fd_sc_hd__inv_2 _4597_ (.A(_2327_),
    .Y(_0406_));
 sky130_fd_sc_hd__inv_2 _4598_ (.A(_2327_),
    .Y(_0407_));
 sky130_fd_sc_hd__buf_2 _4599_ (.A(_2325_),
    .X(_2328_));
 sky130_fd_sc_hd__inv_2 _4600_ (.A(_2328_),
    .Y(_0408_));
 sky130_fd_sc_hd__inv_2 _4601_ (.A(_2328_),
    .Y(_0409_));
 sky130_fd_sc_hd__inv_2 _4602_ (.A(_2328_),
    .Y(_0410_));
 sky130_fd_sc_hd__inv_2 _4603_ (.A(_2328_),
    .Y(_0411_));
 sky130_fd_sc_hd__clkbuf_2 _4604_ (.A(_2325_),
    .X(_2329_));
 sky130_fd_sc_hd__inv_2 _4605_ (.A(_2329_),
    .Y(_0412_));
 sky130_fd_sc_hd__inv_2 _4606_ (.A(_2329_),
    .Y(_0413_));
 sky130_fd_sc_hd__inv_2 _4607_ (.A(_2329_),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_2 _4608_ (.A(_2329_),
    .Y(_0415_));
 sky130_fd_sc_hd__buf_1 _4609_ (.A(_2314_),
    .X(_2330_));
 sky130_fd_sc_hd__clkbuf_2 _4610_ (.A(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__inv_2 _4611_ (.A(_2331_),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_2 _4612_ (.A(_2331_),
    .Y(_0417_));
 sky130_fd_sc_hd__inv_2 _4613_ (.A(_2331_),
    .Y(_0418_));
 sky130_fd_sc_hd__inv_2 _4614_ (.A(_2331_),
    .Y(_0419_));
 sky130_fd_sc_hd__clkbuf_2 _4615_ (.A(_2330_),
    .X(_2332_));
 sky130_fd_sc_hd__inv_2 _4616_ (.A(_2332_),
    .Y(_0420_));
 sky130_fd_sc_hd__inv_2 _4617_ (.A(_2332_),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_2 _4618_ (.A(_2332_),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_2 _4619_ (.A(_2332_),
    .Y(_0423_));
 sky130_fd_sc_hd__clkbuf_2 _4620_ (.A(_2330_),
    .X(_2333_));
 sky130_fd_sc_hd__inv_2 _4621_ (.A(_2333_),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_2 _4622_ (.A(_2333_),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_2 _4623_ (.A(_2333_),
    .Y(_0426_));
 sky130_fd_sc_hd__inv_2 _4624_ (.A(_2333_),
    .Y(_0427_));
 sky130_fd_sc_hd__clkbuf_2 _4625_ (.A(_2330_),
    .X(_2334_));
 sky130_fd_sc_hd__inv_2 _4626_ (.A(_2334_),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _4627_ (.A(_2334_),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_2 _4628_ (.A(_2334_),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _4629_ (.A(_2334_),
    .Y(_0431_));
 sky130_fd_sc_hd__clkbuf_2 _4630_ (.A(_2191_),
    .X(_2335_));
 sky130_fd_sc_hd__buf_1 _4631_ (.A(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__clkbuf_2 _4632_ (.A(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__inv_2 _4633_ (.A(_2337_),
    .Y(_0432_));
 sky130_fd_sc_hd__inv_2 _4634_ (.A(_2337_),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_2 _4635_ (.A(_2337_),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_2 _4636_ (.A(_2337_),
    .Y(_0435_));
 sky130_fd_sc_hd__clkbuf_2 _4637_ (.A(_2336_),
    .X(_2338_));
 sky130_fd_sc_hd__inv_2 _4638_ (.A(_2338_),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_2 _4639_ (.A(_2338_),
    .Y(_0437_));
 sky130_fd_sc_hd__inv_2 _4640_ (.A(_2338_),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_2 _4641_ (.A(_2338_),
    .Y(_0439_));
 sky130_fd_sc_hd__clkbuf_2 _4642_ (.A(_2336_),
    .X(_2339_));
 sky130_fd_sc_hd__inv_2 _4643_ (.A(_2339_),
    .Y(_0440_));
 sky130_fd_sc_hd__inv_2 _4644_ (.A(_2339_),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _4645_ (.A(_2339_),
    .Y(_0442_));
 sky130_fd_sc_hd__inv_2 _4646_ (.A(_2339_),
    .Y(_0443_));
 sky130_fd_sc_hd__clkbuf_2 _4647_ (.A(_2336_),
    .X(_2340_));
 sky130_fd_sc_hd__inv_2 _4648_ (.A(_2340_),
    .Y(_0444_));
 sky130_fd_sc_hd__inv_2 _4649_ (.A(_2340_),
    .Y(_0445_));
 sky130_fd_sc_hd__inv_2 _4650_ (.A(_2340_),
    .Y(_0446_));
 sky130_fd_sc_hd__inv_2 _4651_ (.A(_2340_),
    .Y(_0447_));
 sky130_fd_sc_hd__buf_1 _4652_ (.A(_2335_),
    .X(_2341_));
 sky130_fd_sc_hd__clkbuf_2 _4653_ (.A(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__inv_2 _4654_ (.A(_2342_),
    .Y(_0448_));
 sky130_fd_sc_hd__inv_2 _4655_ (.A(_2342_),
    .Y(_0449_));
 sky130_fd_sc_hd__inv_2 _4656_ (.A(_2342_),
    .Y(_0450_));
 sky130_fd_sc_hd__inv_2 _4657_ (.A(_2342_),
    .Y(_0451_));
 sky130_fd_sc_hd__clkbuf_2 _4658_ (.A(_2341_),
    .X(_2343_));
 sky130_fd_sc_hd__inv_2 _4659_ (.A(_2343_),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _4660_ (.A(_2343_),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_2 _4661_ (.A(_2343_),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _4662_ (.A(_2343_),
    .Y(_0455_));
 sky130_fd_sc_hd__clkbuf_2 _4663_ (.A(_2341_),
    .X(_2344_));
 sky130_fd_sc_hd__inv_2 _4664_ (.A(_2344_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _4665_ (.A(_2344_),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _4666_ (.A(_2344_),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _4667_ (.A(_2344_),
    .Y(_0459_));
 sky130_fd_sc_hd__clkbuf_2 _4668_ (.A(_2341_),
    .X(_2345_));
 sky130_fd_sc_hd__inv_2 _4669_ (.A(_2345_),
    .Y(_0460_));
 sky130_fd_sc_hd__inv_2 _4670_ (.A(_2345_),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_2 _4671_ (.A(_2345_),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_2 _4672_ (.A(_2345_),
    .Y(_0463_));
 sky130_fd_sc_hd__buf_1 _4673_ (.A(_2335_),
    .X(_2346_));
 sky130_fd_sc_hd__clkbuf_2 _4674_ (.A(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__inv_2 _4675_ (.A(_2347_),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_2 _4676_ (.A(_2347_),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _4677_ (.A(_2347_),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_2 _4678_ (.A(_2347_),
    .Y(_0467_));
 sky130_fd_sc_hd__clkbuf_2 _4679_ (.A(_2346_),
    .X(_2348_));
 sky130_fd_sc_hd__inv_2 _4680_ (.A(_2348_),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _4681_ (.A(_2348_),
    .Y(_0469_));
 sky130_fd_sc_hd__inv_2 _4682_ (.A(_2348_),
    .Y(_0470_));
 sky130_fd_sc_hd__inv_2 _4683_ (.A(_2348_),
    .Y(_0471_));
 sky130_fd_sc_hd__clkbuf_2 _4684_ (.A(_2346_),
    .X(_2349_));
 sky130_fd_sc_hd__inv_2 _4685_ (.A(_2349_),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _4686_ (.A(_2349_),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _4687_ (.A(_2349_),
    .Y(_0474_));
 sky130_fd_sc_hd__inv_2 _4688_ (.A(_2349_),
    .Y(_0475_));
 sky130_fd_sc_hd__clkbuf_2 _4689_ (.A(_2346_),
    .X(_2350_));
 sky130_fd_sc_hd__inv_2 _4690_ (.A(_2350_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _4691_ (.A(_2350_),
    .Y(_0477_));
 sky130_fd_sc_hd__inv_2 _4692_ (.A(_2350_),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _4693_ (.A(_2350_),
    .Y(_0479_));
 sky130_fd_sc_hd__buf_1 _4694_ (.A(_2335_),
    .X(_2351_));
 sky130_fd_sc_hd__clkbuf_2 _4695_ (.A(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__inv_2 _4696_ (.A(_2352_),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_2 _4697_ (.A(_2352_),
    .Y(_0481_));
 sky130_fd_sc_hd__inv_2 _4698_ (.A(_2352_),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_2 _4699_ (.A(_2352_),
    .Y(_0483_));
 sky130_fd_sc_hd__clkbuf_2 _4700_ (.A(_2351_),
    .X(_2353_));
 sky130_fd_sc_hd__inv_2 _4701_ (.A(_2353_),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _4702_ (.A(_2353_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _4703_ (.A(_2353_),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_2 _4704_ (.A(_2353_),
    .Y(_0487_));
 sky130_fd_sc_hd__clkbuf_2 _4705_ (.A(_2351_),
    .X(_2354_));
 sky130_fd_sc_hd__inv_2 _4706_ (.A(_2354_),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _4707_ (.A(_2354_),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _4708_ (.A(_2354_),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_2 _4709_ (.A(_2354_),
    .Y(_0491_));
 sky130_fd_sc_hd__clkbuf_2 _4710_ (.A(_2351_),
    .X(_2355_));
 sky130_fd_sc_hd__inv_2 _4711_ (.A(_2355_),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _4712_ (.A(_2355_),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_2 _4713_ (.A(_2355_),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _4714_ (.A(_2355_),
    .Y(_0495_));
 sky130_fd_sc_hd__buf_1 _4715_ (.A(_2192_),
    .X(_2356_));
 sky130_fd_sc_hd__clkbuf_2 _4716_ (.A(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__inv_2 _4717_ (.A(_2357_),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _4718_ (.A(_2357_),
    .Y(_0497_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(_2357_),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _4720_ (.A(_2357_),
    .Y(_0499_));
 sky130_fd_sc_hd__clkbuf_2 _4721_ (.A(_2356_),
    .X(_2358_));
 sky130_fd_sc_hd__inv_2 _4722_ (.A(_2358_),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _4723_ (.A(_2358_),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _4724_ (.A(_2358_),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _4725_ (.A(_2358_),
    .Y(_0503_));
 sky130_fd_sc_hd__clkbuf_2 _4726_ (.A(_2356_),
    .X(_2359_));
 sky130_fd_sc_hd__inv_2 _4727_ (.A(_2359_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _4728_ (.A(_2359_),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _4729_ (.A(_2359_),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _4730_ (.A(_2359_),
    .Y(_0507_));
 sky130_fd_sc_hd__clkbuf_2 _4731_ (.A(_2356_),
    .X(_2360_));
 sky130_fd_sc_hd__inv_2 _4732_ (.A(_2360_),
    .Y(_0508_));
 sky130_fd_sc_hd__inv_2 _4733_ (.A(_2360_),
    .Y(_0509_));
 sky130_fd_sc_hd__inv_2 _4734_ (.A(_2360_),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_2 _4735_ (.A(_2360_),
    .Y(_0511_));
 sky130_fd_sc_hd__buf_1 _4736_ (.A(_2192_),
    .X(_2361_));
 sky130_fd_sc_hd__clkbuf_2 _4737_ (.A(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__inv_2 _4738_ (.A(_2362_),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_2 _4739_ (.A(_2362_),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _4740_ (.A(_2362_),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_2 _4741_ (.A(_2362_),
    .Y(_0515_));
 sky130_fd_sc_hd__clkbuf_2 _4742_ (.A(_2361_),
    .X(_2363_));
 sky130_fd_sc_hd__inv_2 _4743_ (.A(_2363_),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _4744_ (.A(_2363_),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_2 _4745_ (.A(_2363_),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_2 _4746_ (.A(_2363_),
    .Y(_0519_));
 sky130_fd_sc_hd__clkbuf_2 _4747_ (.A(_2361_),
    .X(_2364_));
 sky130_fd_sc_hd__inv_2 _4748_ (.A(_2364_),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _4749_ (.A(_2364_),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _4750_ (.A(_2364_),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _4751_ (.A(_2364_),
    .Y(_0523_));
 sky130_fd_sc_hd__clkbuf_2 _4752_ (.A(_2361_),
    .X(_2365_));
 sky130_fd_sc_hd__inv_2 _4753_ (.A(_2365_),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _4754_ (.A(_2365_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _4755_ (.A(_2365_),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_2 _4756_ (.A(_2365_),
    .Y(_0527_));
 sky130_fd_sc_hd__clkbuf_2 _4757_ (.A(_2197_),
    .X(_2366_));
 sky130_fd_sc_hd__inv_2 _4758_ (.A(_2366_),
    .Y(_0528_));
 sky130_fd_sc_hd__inv_2 _4759_ (.A(_2366_),
    .Y(_0529_));
 sky130_fd_sc_hd__inv_2 _4760_ (.A(_2366_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _4761_ (.A(_2366_),
    .Y(_0531_));
 sky130_fd_sc_hd__clkbuf_2 _4762_ (.A(_2197_),
    .X(_2367_));
 sky130_fd_sc_hd__inv_2 _4763_ (.A(_2367_),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_2 _4764_ (.A(_2367_),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _4765_ (.A(_2367_),
    .Y(_0534_));
 sky130_fd_sc_hd__inv_2 _4766_ (.A(_2367_),
    .Y(_0535_));
 sky130_fd_sc_hd__inv_2 _4767_ (.A(_2193_),
    .Y(_0536_));
 sky130_fd_sc_hd__dfrtp_1 _4768_ (.CLK(clknet_leaf_5_clk),
    .D(_0537_),
    .RESET_B(_0004_),
    .Q(\input_a[14][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4769_ (.CLK(clknet_leaf_4_clk),
    .D(_0538_),
    .RESET_B(_0005_),
    .Q(\output_c[15][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4770_ (.CLK(clknet_leaf_4_clk),
    .D(_0539_),
    .RESET_B(_0006_),
    .Q(\output_c[15][1] ));
 sky130_fd_sc_hd__dfrtp_1 _4771_ (.CLK(clknet_leaf_5_clk),
    .D(_0540_),
    .RESET_B(_0007_),
    .Q(\output_c[15][2] ));
 sky130_fd_sc_hd__dfrtp_1 _4772_ (.CLK(clknet_leaf_5_clk),
    .D(_0541_),
    .RESET_B(_0008_),
    .Q(\output_c[15][3] ));
 sky130_fd_sc_hd__dfrtp_1 _4773_ (.CLK(clknet_leaf_5_clk),
    .D(_0542_),
    .RESET_B(_0009_),
    .Q(\output_c[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _4774_ (.CLK(clknet_leaf_5_clk),
    .D(_0543_),
    .RESET_B(_0010_),
    .Q(\output_c[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _4775_ (.CLK(clknet_leaf_5_clk),
    .D(_0544_),
    .RESET_B(_0011_),
    .Q(\output_c[15][6] ));
 sky130_fd_sc_hd__dfrtp_1 _4776_ (.CLK(clknet_leaf_5_clk),
    .D(_0545_),
    .RESET_B(_0012_),
    .Q(\output_c[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _4777_ (.CLK(clknet_leaf_6_clk),
    .D(_0546_),
    .RESET_B(_0013_),
    .Q(\output_c[15][8] ));
 sky130_fd_sc_hd__dfrtp_1 _4778_ (.CLK(clknet_leaf_5_clk),
    .D(_0547_),
    .RESET_B(_0014_),
    .Q(\output_c[15][9] ));
 sky130_fd_sc_hd__dfrtp_1 _4779_ (.CLK(clknet_leaf_6_clk),
    .D(_0548_),
    .RESET_B(_0015_),
    .Q(\output_c[15][10] ));
 sky130_fd_sc_hd__dfrtp_1 _4780_ (.CLK(clknet_leaf_7_clk),
    .D(_0549_),
    .RESET_B(_0016_),
    .Q(\output_c[15][11] ));
 sky130_fd_sc_hd__dfrtp_1 _4781_ (.CLK(clknet_leaf_7_clk),
    .D(_0550_),
    .RESET_B(_0017_),
    .Q(\output_c[15][12] ));
 sky130_fd_sc_hd__dfrtp_1 _4782_ (.CLK(clknet_leaf_7_clk),
    .D(_0551_),
    .RESET_B(_0018_),
    .Q(\output_c[15][13] ));
 sky130_fd_sc_hd__dfrtp_1 _4783_ (.CLK(clknet_leaf_7_clk),
    .D(_0552_),
    .RESET_B(_0019_),
    .Q(\output_c[15][14] ));
 sky130_fd_sc_hd__dfrtp_1 _4784_ (.CLK(clknet_leaf_7_clk),
    .D(_0553_),
    .RESET_B(_0020_),
    .Q(\output_c[15][15] ));
 sky130_fd_sc_hd__dfrtp_1 _4785_ (.CLK(clknet_leaf_7_clk),
    .D(_0554_),
    .RESET_B(_0021_),
    .Q(\output_c[15][16] ));
 sky130_fd_sc_hd__dfrtp_1 _4786_ (.CLK(clknet_leaf_7_clk),
    .D(_0555_),
    .RESET_B(_0022_),
    .Q(\output_c[15][17] ));
 sky130_fd_sc_hd__dfrtp_1 _4787_ (.CLK(clknet_leaf_7_clk),
    .D(_0556_),
    .RESET_B(_0023_),
    .Q(\output_c[15][18] ));
 sky130_fd_sc_hd__dfrtp_1 _4788_ (.CLK(clknet_leaf_7_clk),
    .D(_0557_),
    .RESET_B(_0024_),
    .Q(\output_c[15][19] ));
 sky130_fd_sc_hd__dfrtp_1 _4789_ (.CLK(clknet_leaf_7_clk),
    .D(_0558_),
    .RESET_B(_0025_),
    .Q(\output_c[15][20] ));
 sky130_fd_sc_hd__dfrtp_1 _4790_ (.CLK(clknet_leaf_7_clk),
    .D(_0559_),
    .RESET_B(_0026_),
    .Q(\output_c[15][21] ));
 sky130_fd_sc_hd__dfrtp_1 _4791_ (.CLK(clknet_leaf_8_clk),
    .D(net145),
    .RESET_B(_0027_),
    .Q(\output_c[15][22] ));
 sky130_fd_sc_hd__dfrtp_1 _4792_ (.CLK(clknet_leaf_8_clk),
    .D(_0561_),
    .RESET_B(_0028_),
    .Q(\output_c[15][23] ));
 sky130_fd_sc_hd__dfrtp_1 _4793_ (.CLK(clknet_leaf_8_clk),
    .D(_0562_),
    .RESET_B(_0029_),
    .Q(\output_c[15][24] ));
 sky130_fd_sc_hd__dfrtp_1 _4794_ (.CLK(clknet_leaf_8_clk),
    .D(_0563_),
    .RESET_B(_0030_),
    .Q(\output_c[15][25] ));
 sky130_fd_sc_hd__dfrtp_1 _4795_ (.CLK(clknet_leaf_8_clk),
    .D(_0564_),
    .RESET_B(_0031_),
    .Q(\output_c[15][26] ));
 sky130_fd_sc_hd__dfrtp_1 _4796_ (.CLK(clknet_leaf_5_clk),
    .D(_0565_),
    .RESET_B(_0032_),
    .Q(\output_c[15][27] ));
 sky130_fd_sc_hd__dfrtp_1 _4797_ (.CLK(clknet_leaf_5_clk),
    .D(_0566_),
    .RESET_B(_0033_),
    .Q(\output_c[15][28] ));
 sky130_fd_sc_hd__dfrtp_1 _4798_ (.CLK(clknet_leaf_5_clk),
    .D(_0567_),
    .RESET_B(_0034_),
    .Q(\output_c[15][29] ));
 sky130_fd_sc_hd__dfrtp_1 _4799_ (.CLK(clknet_leaf_5_clk),
    .D(_0568_),
    .RESET_B(_0035_),
    .Q(\output_c[15][30] ));
 sky130_fd_sc_hd__dfrtp_1 _4800_ (.CLK(clknet_leaf_5_clk),
    .D(_0569_),
    .RESET_B(_0036_),
    .Q(\output_c[15][31] ));
 sky130_fd_sc_hd__dfrtp_1 _4801_ (.CLK(clknet_leaf_4_clk),
    .D(_0000_),
    .RESET_B(_0037_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4802_ (.CLK(clknet_leaf_4_clk),
    .D(_0001_),
    .RESET_B(_0038_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4803_ (.CLK(clknet_leaf_4_clk),
    .D(_0002_),
    .RESET_B(_0039_),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4804_ (.CLK(clknet_leaf_4_clk),
    .D(_0003_),
    .RESET_B(_0040_),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4805_ (.CLK(clknet_leaf_4_clk),
    .D(_0570_),
    .RESET_B(_0041_),
    .Q(\input_a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4806_ (.CLK(clknet_leaf_15_clk),
    .D(_0571_),
    .RESET_B(_0042_),
    .Q(\input_a[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4807_ (.CLK(clknet_leaf_15_clk),
    .D(_0572_),
    .RESET_B(_0043_),
    .Q(\input_a[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4808_ (.CLK(clknet_leaf_26_clk),
    .D(_0573_),
    .RESET_B(_0044_),
    .Q(\input_a[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4809_ (.CLK(clknet_leaf_26_clk),
    .D(_0574_),
    .RESET_B(_0045_),
    .Q(\input_a[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4810_ (.CLK(clknet_leaf_36_clk),
    .D(_0575_),
    .RESET_B(_0046_),
    .Q(\input_a[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4811_ (.CLK(clknet_leaf_36_clk),
    .D(_0576_),
    .RESET_B(_0047_),
    .Q(\input_a[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4812_ (.CLK(clknet_leaf_4_clk),
    .D(_0577_),
    .RESET_B(_0048_),
    .Q(\input_a[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4813_ (.CLK(clknet_leaf_4_clk),
    .D(_0578_),
    .RESET_B(_0049_),
    .Q(\input_a[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4814_ (.CLK(clknet_leaf_4_clk),
    .D(_0579_),
    .RESET_B(_0050_),
    .Q(\input_a[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4815_ (.CLK(clknet_leaf_4_clk),
    .D(_0580_),
    .RESET_B(_0051_),
    .Q(\input_a[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4816_ (.CLK(clknet_leaf_15_clk),
    .D(_0581_),
    .RESET_B(_0052_),
    .Q(\input_a[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4817_ (.CLK(clknet_leaf_15_clk),
    .D(_0582_),
    .RESET_B(_0053_),
    .Q(\input_a[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4818_ (.CLK(clknet_leaf_15_clk),
    .D(_0583_),
    .RESET_B(_0054_),
    .Q(\input_a[12][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4819_ (.CLK(clknet_leaf_15_clk),
    .D(_0584_),
    .RESET_B(_0055_),
    .Q(\input_a[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4820_ (.CLK(clknet_leaf_15_clk),
    .D(_0585_),
    .RESET_B(_0056_),
    .Q(\input_b[15][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4821_ (.CLK(clknet_leaf_15_clk),
    .D(_0586_),
    .RESET_B(_0057_),
    .Q(\output_c[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4822_ (.CLK(clknet_leaf_15_clk),
    .D(_0587_),
    .RESET_B(_0058_),
    .Q(\output_c[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _4823_ (.CLK(clknet_leaf_15_clk),
    .D(net414),
    .RESET_B(_0059_),
    .Q(\output_c[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _4824_ (.CLK(clknet_leaf_15_clk),
    .D(_0589_),
    .RESET_B(_0060_),
    .Q(\output_c[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _4825_ (.CLK(clknet_leaf_15_clk),
    .D(_0590_),
    .RESET_B(_0061_),
    .Q(\output_c[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _4826_ (.CLK(clknet_leaf_15_clk),
    .D(_0591_),
    .RESET_B(_0062_),
    .Q(\output_c[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _4827_ (.CLK(clknet_leaf_14_clk),
    .D(_0592_),
    .RESET_B(_0063_),
    .Q(\output_c[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _4828_ (.CLK(clknet_leaf_14_clk),
    .D(_0593_),
    .RESET_B(_0064_),
    .Q(\output_c[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _4829_ (.CLK(clknet_leaf_13_clk),
    .D(_0594_),
    .RESET_B(_0065_),
    .Q(\output_c[0][8] ));
 sky130_fd_sc_hd__dfrtp_1 _4830_ (.CLK(clknet_leaf_13_clk),
    .D(_0595_),
    .RESET_B(_0066_),
    .Q(\output_c[0][9] ));
 sky130_fd_sc_hd__dfrtp_1 _4831_ (.CLK(clknet_leaf_13_clk),
    .D(_0596_),
    .RESET_B(_0067_),
    .Q(\output_c[0][10] ));
 sky130_fd_sc_hd__dfrtp_1 _4832_ (.CLK(clknet_leaf_13_clk),
    .D(_0597_),
    .RESET_B(_0068_),
    .Q(\output_c[0][11] ));
 sky130_fd_sc_hd__dfrtp_1 _4833_ (.CLK(clknet_leaf_13_clk),
    .D(_0598_),
    .RESET_B(_0069_),
    .Q(\output_c[0][12] ));
 sky130_fd_sc_hd__dfrtp_1 _4834_ (.CLK(clknet_leaf_13_clk),
    .D(_0599_),
    .RESET_B(_0070_),
    .Q(\output_c[0][13] ));
 sky130_fd_sc_hd__dfrtp_1 _4835_ (.CLK(clknet_leaf_13_clk),
    .D(_0600_),
    .RESET_B(_0071_),
    .Q(\output_c[0][14] ));
 sky130_fd_sc_hd__dfrtp_1 _4836_ (.CLK(clknet_leaf_13_clk),
    .D(_0601_),
    .RESET_B(_0072_),
    .Q(\output_c[0][15] ));
 sky130_fd_sc_hd__dfrtp_1 _4837_ (.CLK(clknet_leaf_13_clk),
    .D(_0602_),
    .RESET_B(_0073_),
    .Q(\output_c[0][16] ));
 sky130_fd_sc_hd__dfrtp_1 _4838_ (.CLK(clknet_leaf_13_clk),
    .D(_0603_),
    .RESET_B(_0074_),
    .Q(\output_c[0][17] ));
 sky130_fd_sc_hd__dfrtp_1 _4839_ (.CLK(clknet_leaf_13_clk),
    .D(_0604_),
    .RESET_B(_0075_),
    .Q(\output_c[0][18] ));
 sky130_fd_sc_hd__dfrtp_1 _4840_ (.CLK(clknet_leaf_13_clk),
    .D(_0605_),
    .RESET_B(_0076_),
    .Q(\output_c[0][19] ));
 sky130_fd_sc_hd__dfrtp_1 _4841_ (.CLK(clknet_leaf_17_clk),
    .D(_0606_),
    .RESET_B(_0077_),
    .Q(\output_c[0][20] ));
 sky130_fd_sc_hd__dfrtp_1 _4842_ (.CLK(clknet_leaf_17_clk),
    .D(_0607_),
    .RESET_B(_0078_),
    .Q(\output_c[0][21] ));
 sky130_fd_sc_hd__dfrtp_1 _4843_ (.CLK(clknet_leaf_17_clk),
    .D(_0608_),
    .RESET_B(_0079_),
    .Q(\output_c[0][22] ));
 sky130_fd_sc_hd__dfrtp_1 _4844_ (.CLK(clknet_leaf_17_clk),
    .D(_0609_),
    .RESET_B(_0080_),
    .Q(\output_c[0][23] ));
 sky130_fd_sc_hd__dfrtp_1 _4845_ (.CLK(clknet_leaf_16_clk),
    .D(_0610_),
    .RESET_B(_0081_),
    .Q(\output_c[0][24] ));
 sky130_fd_sc_hd__dfrtp_1 _4846_ (.CLK(clknet_leaf_16_clk),
    .D(_0611_),
    .RESET_B(_0082_),
    .Q(\output_c[0][25] ));
 sky130_fd_sc_hd__dfrtp_1 _4847_ (.CLK(clknet_leaf_16_clk),
    .D(_0612_),
    .RESET_B(_0083_),
    .Q(\output_c[0][26] ));
 sky130_fd_sc_hd__dfrtp_1 _4848_ (.CLK(clknet_leaf_17_clk),
    .D(_0613_),
    .RESET_B(_0084_),
    .Q(\output_c[0][27] ));
 sky130_fd_sc_hd__dfrtp_1 _4849_ (.CLK(clknet_leaf_16_clk),
    .D(_0614_),
    .RESET_B(_0085_),
    .Q(\output_c[0][28] ));
 sky130_fd_sc_hd__dfrtp_1 _4850_ (.CLK(clknet_leaf_16_clk),
    .D(_0615_),
    .RESET_B(_0086_),
    .Q(\output_c[0][29] ));
 sky130_fd_sc_hd__dfrtp_1 _4851_ (.CLK(clknet_leaf_16_clk),
    .D(_0616_),
    .RESET_B(_0087_),
    .Q(\output_c[0][30] ));
 sky130_fd_sc_hd__dfrtp_1 _4852_ (.CLK(clknet_leaf_16_clk),
    .D(_0617_),
    .RESET_B(_0088_),
    .Q(\output_c[0][31] ));
 sky130_fd_sc_hd__dfrtp_1 _4853_ (.CLK(clknet_leaf_15_clk),
    .D(_0618_),
    .RESET_B(_0089_),
    .Q(\output_c[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4854_ (.CLK(clknet_leaf_26_clk),
    .D(_0619_),
    .RESET_B(_0090_),
    .Q(\output_c[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _4855_ (.CLK(clknet_leaf_15_clk),
    .D(net443),
    .RESET_B(_0091_),
    .Q(\output_c[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _4856_ (.CLK(clknet_leaf_25_clk),
    .D(_0621_),
    .RESET_B(_0092_),
    .Q(\output_c[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _4857_ (.CLK(clknet_leaf_25_clk),
    .D(_0622_),
    .RESET_B(_0093_),
    .Q(\output_c[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _4858_ (.CLK(clknet_leaf_16_clk),
    .D(_0623_),
    .RESET_B(_0094_),
    .Q(\output_c[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _4859_ (.CLK(clknet_leaf_25_clk),
    .D(_0624_),
    .RESET_B(_0095_),
    .Q(\output_c[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _4860_ (.CLK(clknet_leaf_16_clk),
    .D(_0625_),
    .RESET_B(_0096_),
    .Q(\output_c[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _4861_ (.CLK(clknet_leaf_16_clk),
    .D(_0626_),
    .RESET_B(_0097_),
    .Q(\output_c[1][8] ));
 sky130_fd_sc_hd__dfrtp_1 _4862_ (.CLK(clknet_leaf_16_clk),
    .D(_0627_),
    .RESET_B(_0098_),
    .Q(\output_c[1][9] ));
 sky130_fd_sc_hd__dfrtp_1 _4863_ (.CLK(clknet_leaf_16_clk),
    .D(_0628_),
    .RESET_B(_0099_),
    .Q(\output_c[1][10] ));
 sky130_fd_sc_hd__dfrtp_1 _4864_ (.CLK(clknet_leaf_16_clk),
    .D(_0629_),
    .RESET_B(_0100_),
    .Q(\output_c[1][11] ));
 sky130_fd_sc_hd__dfrtp_1 _4865_ (.CLK(clknet_leaf_16_clk),
    .D(_0630_),
    .RESET_B(_0101_),
    .Q(\output_c[1][12] ));
 sky130_fd_sc_hd__dfrtp_1 _4866_ (.CLK(clknet_leaf_16_clk),
    .D(_0631_),
    .RESET_B(_0102_),
    .Q(\output_c[1][13] ));
 sky130_fd_sc_hd__dfrtp_1 _4867_ (.CLK(clknet_leaf_16_clk),
    .D(_0632_),
    .RESET_B(_0103_),
    .Q(\output_c[1][14] ));
 sky130_fd_sc_hd__dfrtp_1 _4868_ (.CLK(clknet_leaf_19_clk),
    .D(_0633_),
    .RESET_B(_0104_),
    .Q(\output_c[1][15] ));
 sky130_fd_sc_hd__dfrtp_1 _4869_ (.CLK(clknet_leaf_22_clk),
    .D(_0634_),
    .RESET_B(_0105_),
    .Q(\output_c[1][16] ));
 sky130_fd_sc_hd__dfrtp_1 _4870_ (.CLK(clknet_leaf_19_clk),
    .D(_0635_),
    .RESET_B(_0106_),
    .Q(\output_c[1][17] ));
 sky130_fd_sc_hd__dfrtp_1 _4871_ (.CLK(clknet_leaf_19_clk),
    .D(_0636_),
    .RESET_B(_0107_),
    .Q(\output_c[1][18] ));
 sky130_fd_sc_hd__dfrtp_1 _4872_ (.CLK(clknet_leaf_21_clk),
    .D(_0637_),
    .RESET_B(_0108_),
    .Q(\output_c[1][19] ));
 sky130_fd_sc_hd__dfrtp_1 _4873_ (.CLK(clknet_leaf_22_clk),
    .D(_0638_),
    .RESET_B(_0109_),
    .Q(\output_c[1][20] ));
 sky130_fd_sc_hd__dfrtp_1 _4874_ (.CLK(clknet_leaf_22_clk),
    .D(_0639_),
    .RESET_B(_0110_),
    .Q(\output_c[1][21] ));
 sky130_fd_sc_hd__dfrtp_1 _4875_ (.CLK(clknet_leaf_22_clk),
    .D(_0640_),
    .RESET_B(_0111_),
    .Q(\output_c[1][22] ));
 sky130_fd_sc_hd__dfrtp_1 _4876_ (.CLK(clknet_leaf_25_clk),
    .D(_0641_),
    .RESET_B(_0112_),
    .Q(\output_c[1][23] ));
 sky130_fd_sc_hd__dfrtp_1 _4877_ (.CLK(clknet_leaf_25_clk),
    .D(_0642_),
    .RESET_B(_0113_),
    .Q(\output_c[1][24] ));
 sky130_fd_sc_hd__dfrtp_1 _4878_ (.CLK(clknet_leaf_25_clk),
    .D(_0643_),
    .RESET_B(_0114_),
    .Q(\output_c[1][25] ));
 sky130_fd_sc_hd__dfrtp_1 _4879_ (.CLK(clknet_leaf_24_clk),
    .D(_0644_),
    .RESET_B(_0115_),
    .Q(\output_c[1][26] ));
 sky130_fd_sc_hd__dfrtp_1 _4880_ (.CLK(clknet_leaf_24_clk),
    .D(_0645_),
    .RESET_B(_0116_),
    .Q(\output_c[1][27] ));
 sky130_fd_sc_hd__dfrtp_1 _4881_ (.CLK(clknet_leaf_24_clk),
    .D(_0646_),
    .RESET_B(_0117_),
    .Q(\output_c[1][28] ));
 sky130_fd_sc_hd__dfrtp_1 _4882_ (.CLK(clknet_leaf_24_clk),
    .D(_0647_),
    .RESET_B(_0118_),
    .Q(\output_c[1][29] ));
 sky130_fd_sc_hd__dfrtp_1 _4883_ (.CLK(clknet_leaf_25_clk),
    .D(_0648_),
    .RESET_B(_0119_),
    .Q(\output_c[1][30] ));
 sky130_fd_sc_hd__dfrtp_1 _4884_ (.CLK(clknet_leaf_25_clk),
    .D(_0649_),
    .RESET_B(_0120_),
    .Q(\output_c[1][31] ));
 sky130_fd_sc_hd__dfrtp_1 _4885_ (.CLK(clknet_leaf_26_clk),
    .D(_0650_),
    .RESET_B(_0121_),
    .Q(\output_c[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4886_ (.CLK(clknet_leaf_26_clk),
    .D(_0651_),
    .RESET_B(_0122_),
    .Q(\output_c[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _4887_ (.CLK(clknet_leaf_25_clk),
    .D(net351),
    .RESET_B(_0123_),
    .Q(\output_c[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _4888_ (.CLK(clknet_leaf_25_clk),
    .D(_0653_),
    .RESET_B(_0124_),
    .Q(\output_c[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _4889_ (.CLK(clknet_leaf_24_clk),
    .D(_0654_),
    .RESET_B(_0125_),
    .Q(\output_c[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _4890_ (.CLK(clknet_leaf_24_clk),
    .D(_0655_),
    .RESET_B(_0126_),
    .Q(\output_c[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _4891_ (.CLK(clknet_leaf_24_clk),
    .D(_0656_),
    .RESET_B(_0127_),
    .Q(\output_c[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _4892_ (.CLK(clknet_leaf_24_clk),
    .D(_0657_),
    .RESET_B(_0128_),
    .Q(\output_c[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _4893_ (.CLK(clknet_leaf_23_clk),
    .D(_0658_),
    .RESET_B(_0129_),
    .Q(\output_c[2][8] ));
 sky130_fd_sc_hd__dfrtp_1 _4894_ (.CLK(clknet_leaf_23_clk),
    .D(_0659_),
    .RESET_B(_0130_),
    .Q(\output_c[2][9] ));
 sky130_fd_sc_hd__dfrtp_1 _4895_ (.CLK(clknet_leaf_23_clk),
    .D(_0660_),
    .RESET_B(_0131_),
    .Q(\output_c[2][10] ));
 sky130_fd_sc_hd__dfrtp_1 _4896_ (.CLK(clknet_leaf_23_clk),
    .D(_0661_),
    .RESET_B(_0132_),
    .Q(\output_c[2][11] ));
 sky130_fd_sc_hd__dfrtp_1 _4897_ (.CLK(clknet_leaf_23_clk),
    .D(_0662_),
    .RESET_B(_0133_),
    .Q(\output_c[2][12] ));
 sky130_fd_sc_hd__dfrtp_1 _4898_ (.CLK(clknet_leaf_23_clk),
    .D(_0663_),
    .RESET_B(_0134_),
    .Q(\output_c[2][13] ));
 sky130_fd_sc_hd__dfrtp_1 _4899_ (.CLK(clknet_leaf_23_clk),
    .D(_0664_),
    .RESET_B(_0135_),
    .Q(\output_c[2][14] ));
 sky130_fd_sc_hd__dfrtp_1 _4900_ (.CLK(clknet_leaf_24_clk),
    .D(_0665_),
    .RESET_B(_0136_),
    .Q(\output_c[2][15] ));
 sky130_fd_sc_hd__dfrtp_1 _4901_ (.CLK(clknet_leaf_28_clk),
    .D(_0666_),
    .RESET_B(_0137_),
    .Q(\output_c[2][16] ));
 sky130_fd_sc_hd__dfrtp_1 _4902_ (.CLK(clknet_leaf_28_clk),
    .D(_0667_),
    .RESET_B(_0138_),
    .Q(\output_c[2][17] ));
 sky130_fd_sc_hd__dfrtp_1 _4903_ (.CLK(clknet_leaf_28_clk),
    .D(_0668_),
    .RESET_B(_0139_),
    .Q(\output_c[2][18] ));
 sky130_fd_sc_hd__dfrtp_1 _4904_ (.CLK(clknet_leaf_28_clk),
    .D(_0669_),
    .RESET_B(_0140_),
    .Q(\output_c[2][19] ));
 sky130_fd_sc_hd__dfrtp_1 _4905_ (.CLK(clknet_leaf_28_clk),
    .D(_0670_),
    .RESET_B(_0141_),
    .Q(\output_c[2][20] ));
 sky130_fd_sc_hd__dfrtp_1 _4906_ (.CLK(clknet_leaf_28_clk),
    .D(_0671_),
    .RESET_B(_0142_),
    .Q(\output_c[2][21] ));
 sky130_fd_sc_hd__dfrtp_1 _4907_ (.CLK(clknet_leaf_28_clk),
    .D(_0672_),
    .RESET_B(_0143_),
    .Q(\output_c[2][22] ));
 sky130_fd_sc_hd__dfrtp_1 _4908_ (.CLK(clknet_leaf_28_clk),
    .D(_0673_),
    .RESET_B(_0144_),
    .Q(\output_c[2][23] ));
 sky130_fd_sc_hd__dfrtp_1 _4909_ (.CLK(clknet_leaf_28_clk),
    .D(_0674_),
    .RESET_B(_0145_),
    .Q(\output_c[2][24] ));
 sky130_fd_sc_hd__dfrtp_1 _4910_ (.CLK(clknet_leaf_27_clk),
    .D(_0675_),
    .RESET_B(_0146_),
    .Q(\output_c[2][25] ));
 sky130_fd_sc_hd__dfrtp_1 _4911_ (.CLK(clknet_leaf_27_clk),
    .D(_0676_),
    .RESET_B(_0147_),
    .Q(\output_c[2][26] ));
 sky130_fd_sc_hd__dfrtp_1 _4912_ (.CLK(clknet_leaf_28_clk),
    .D(_0677_),
    .RESET_B(_0148_),
    .Q(\output_c[2][27] ));
 sky130_fd_sc_hd__dfrtp_1 _4913_ (.CLK(clknet_leaf_28_clk),
    .D(_0678_),
    .RESET_B(_0149_),
    .Q(\output_c[2][28] ));
 sky130_fd_sc_hd__dfrtp_1 _4914_ (.CLK(clknet_leaf_27_clk),
    .D(_0679_),
    .RESET_B(_0150_),
    .Q(\output_c[2][29] ));
 sky130_fd_sc_hd__dfrtp_1 _4915_ (.CLK(clknet_leaf_26_clk),
    .D(_0680_),
    .RESET_B(_0151_),
    .Q(\output_c[2][30] ));
 sky130_fd_sc_hd__dfrtp_1 _4916_ (.CLK(clknet_leaf_26_clk),
    .D(_0681_),
    .RESET_B(_0152_),
    .Q(\output_c[2][31] ));
 sky130_fd_sc_hd__dfrtp_1 _4917_ (.CLK(clknet_leaf_26_clk),
    .D(_0682_),
    .RESET_B(_0153_),
    .Q(\output_c[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4918_ (.CLK(clknet_leaf_27_clk),
    .D(_0683_),
    .RESET_B(_0154_),
    .Q(\output_c[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _4919_ (.CLK(clknet_leaf_27_clk),
    .D(_0684_),
    .RESET_B(_0155_),
    .Q(\output_c[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _4920_ (.CLK(clknet_leaf_27_clk),
    .D(_0685_),
    .RESET_B(_0156_),
    .Q(\output_c[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _4921_ (.CLK(clknet_leaf_27_clk),
    .D(_0686_),
    .RESET_B(_0157_),
    .Q(\output_c[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _4922_ (.CLK(clknet_leaf_27_clk),
    .D(_0687_),
    .RESET_B(_0158_),
    .Q(\output_c[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _4923_ (.CLK(clknet_leaf_27_clk),
    .D(_0688_),
    .RESET_B(_0159_),
    .Q(\output_c[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _4924_ (.CLK(clknet_leaf_28_clk),
    .D(_0689_),
    .RESET_B(_0160_),
    .Q(\output_c[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _4925_ (.CLK(clknet_leaf_29_clk),
    .D(_0690_),
    .RESET_B(_0161_),
    .Q(\output_c[3][8] ));
 sky130_fd_sc_hd__dfrtp_1 _4926_ (.CLK(clknet_leaf_28_clk),
    .D(_0691_),
    .RESET_B(_0162_),
    .Q(\output_c[3][9] ));
 sky130_fd_sc_hd__dfrtp_1 _4927_ (.CLK(clknet_leaf_29_clk),
    .D(_0692_),
    .RESET_B(_0163_),
    .Q(\output_c[3][10] ));
 sky130_fd_sc_hd__dfrtp_1 _4928_ (.CLK(clknet_leaf_28_clk),
    .D(_0693_),
    .RESET_B(_0164_),
    .Q(\output_c[3][11] ));
 sky130_fd_sc_hd__dfrtp_1 _4929_ (.CLK(clknet_leaf_29_clk),
    .D(_0694_),
    .RESET_B(_0165_),
    .Q(\output_c[3][12] ));
 sky130_fd_sc_hd__dfrtp_1 _4930_ (.CLK(clknet_leaf_29_clk),
    .D(_0695_),
    .RESET_B(_0166_),
    .Q(\output_c[3][13] ));
 sky130_fd_sc_hd__dfrtp_1 _4931_ (.CLK(clknet_leaf_29_clk),
    .D(_0696_),
    .RESET_B(_0167_),
    .Q(\output_c[3][14] ));
 sky130_fd_sc_hd__dfrtp_1 _4932_ (.CLK(clknet_leaf_29_clk),
    .D(_0697_),
    .RESET_B(_0168_),
    .Q(\output_c[3][15] ));
 sky130_fd_sc_hd__dfrtp_1 _4933_ (.CLK(clknet_leaf_29_clk),
    .D(_0698_),
    .RESET_B(_0169_),
    .Q(\output_c[3][16] ));
 sky130_fd_sc_hd__dfrtp_1 _4934_ (.CLK(clknet_leaf_30_clk),
    .D(_0699_),
    .RESET_B(_0170_),
    .Q(\output_c[3][17] ));
 sky130_fd_sc_hd__dfrtp_1 _4935_ (.CLK(clknet_leaf_30_clk),
    .D(_0700_),
    .RESET_B(_0171_),
    .Q(\output_c[3][18] ));
 sky130_fd_sc_hd__dfrtp_1 _4936_ (.CLK(clknet_leaf_30_clk),
    .D(_0701_),
    .RESET_B(_0172_),
    .Q(\output_c[3][19] ));
 sky130_fd_sc_hd__dfrtp_1 _4937_ (.CLK(clknet_leaf_30_clk),
    .D(_0702_),
    .RESET_B(_0173_),
    .Q(\output_c[3][20] ));
 sky130_fd_sc_hd__dfrtp_1 _4938_ (.CLK(clknet_leaf_30_clk),
    .D(_0703_),
    .RESET_B(_0174_),
    .Q(\output_c[3][21] ));
 sky130_fd_sc_hd__dfrtp_1 _4939_ (.CLK(clknet_leaf_29_clk),
    .D(_0704_),
    .RESET_B(_0175_),
    .Q(\output_c[3][22] ));
 sky130_fd_sc_hd__dfrtp_1 _4940_ (.CLK(clknet_leaf_30_clk),
    .D(_0705_),
    .RESET_B(_0176_),
    .Q(\output_c[3][23] ));
 sky130_fd_sc_hd__dfrtp_1 _4941_ (.CLK(clknet_leaf_30_clk),
    .D(_0706_),
    .RESET_B(_0177_),
    .Q(\output_c[3][24] ));
 sky130_fd_sc_hd__dfrtp_1 _4942_ (.CLK(clknet_leaf_31_clk),
    .D(_0707_),
    .RESET_B(_0178_),
    .Q(\output_c[3][25] ));
 sky130_fd_sc_hd__dfrtp_1 _4943_ (.CLK(clknet_leaf_31_clk),
    .D(_0708_),
    .RESET_B(_0179_),
    .Q(\output_c[3][26] ));
 sky130_fd_sc_hd__dfrtp_1 _4944_ (.CLK(clknet_leaf_30_clk),
    .D(_0709_),
    .RESET_B(_0180_),
    .Q(\output_c[3][27] ));
 sky130_fd_sc_hd__dfrtp_1 _4945_ (.CLK(clknet_leaf_29_clk),
    .D(_0710_),
    .RESET_B(_0181_),
    .Q(\output_c[3][28] ));
 sky130_fd_sc_hd__dfrtp_1 _4946_ (.CLK(clknet_leaf_30_clk),
    .D(_0711_),
    .RESET_B(_0182_),
    .Q(\output_c[3][29] ));
 sky130_fd_sc_hd__dfrtp_1 _4947_ (.CLK(clknet_leaf_27_clk),
    .D(net86),
    .RESET_B(_0183_),
    .Q(\output_c[3][30] ));
 sky130_fd_sc_hd__dfrtp_1 _4948_ (.CLK(clknet_leaf_27_clk),
    .D(net46),
    .RESET_B(_0184_),
    .Q(\output_c[3][31] ));
 sky130_fd_sc_hd__dfrtp_1 _4949_ (.CLK(clknet_leaf_36_clk),
    .D(_0714_),
    .RESET_B(_0185_),
    .Q(\output_c[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4950_ (.CLK(clknet_leaf_35_clk),
    .D(_0715_),
    .RESET_B(_0186_),
    .Q(\output_c[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _4951_ (.CLK(clknet_leaf_27_clk),
    .D(net439),
    .RESET_B(_0187_),
    .Q(\output_c[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _4952_ (.CLK(clknet_leaf_27_clk),
    .D(_0717_),
    .RESET_B(_0188_),
    .Q(\output_c[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _4953_ (.CLK(clknet_leaf_32_clk),
    .D(_0718_),
    .RESET_B(_0189_),
    .Q(\output_c[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _4954_ (.CLK(clknet_leaf_32_clk),
    .D(_0719_),
    .RESET_B(_0190_),
    .Q(\output_c[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _4955_ (.CLK(clknet_leaf_32_clk),
    .D(_0720_),
    .RESET_B(_0191_),
    .Q(\output_c[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _4956_ (.CLK(clknet_leaf_32_clk),
    .D(_0721_),
    .RESET_B(_0192_),
    .Q(\output_c[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _4957_ (.CLK(clknet_leaf_31_clk),
    .D(_0722_),
    .RESET_B(_0193_),
    .Q(\output_c[4][8] ));
 sky130_fd_sc_hd__dfrtp_1 _4958_ (.CLK(clknet_leaf_31_clk),
    .D(_0723_),
    .RESET_B(_0194_),
    .Q(\output_c[4][9] ));
 sky130_fd_sc_hd__dfrtp_1 _4959_ (.CLK(clknet_leaf_31_clk),
    .D(_0724_),
    .RESET_B(_0195_),
    .Q(\output_c[4][10] ));
 sky130_fd_sc_hd__dfrtp_1 _4960_ (.CLK(clknet_leaf_31_clk),
    .D(_0725_),
    .RESET_B(_0196_),
    .Q(\output_c[4][11] ));
 sky130_fd_sc_hd__dfrtp_1 _4961_ (.CLK(clknet_leaf_31_clk),
    .D(_0726_),
    .RESET_B(_0197_),
    .Q(\output_c[4][12] ));
 sky130_fd_sc_hd__dfrtp_1 _4962_ (.CLK(clknet_leaf_31_clk),
    .D(_0727_),
    .RESET_B(_0198_),
    .Q(\output_c[4][13] ));
 sky130_fd_sc_hd__dfrtp_1 _4963_ (.CLK(clknet_leaf_31_clk),
    .D(_0728_),
    .RESET_B(_0199_),
    .Q(\output_c[4][14] ));
 sky130_fd_sc_hd__dfrtp_1 _4964_ (.CLK(clknet_leaf_31_clk),
    .D(_0729_),
    .RESET_B(_0200_),
    .Q(\output_c[4][15] ));
 sky130_fd_sc_hd__dfrtp_1 _4965_ (.CLK(clknet_leaf_31_clk),
    .D(_0730_),
    .RESET_B(_0201_),
    .Q(\output_c[4][16] ));
 sky130_fd_sc_hd__dfrtp_1 _4966_ (.CLK(clknet_leaf_31_clk),
    .D(_0731_),
    .RESET_B(_0202_),
    .Q(\output_c[4][17] ));
 sky130_fd_sc_hd__dfrtp_1 _4967_ (.CLK(clknet_leaf_31_clk),
    .D(_0732_),
    .RESET_B(_0203_),
    .Q(\output_c[4][18] ));
 sky130_fd_sc_hd__dfrtp_1 _4968_ (.CLK(clknet_leaf_32_clk),
    .D(_0733_),
    .RESET_B(_0204_),
    .Q(\output_c[4][19] ));
 sky130_fd_sc_hd__dfrtp_1 _4969_ (.CLK(clknet_leaf_33_clk),
    .D(_0734_),
    .RESET_B(_0205_),
    .Q(\output_c[4][20] ));
 sky130_fd_sc_hd__dfrtp_1 _4970_ (.CLK(clknet_leaf_32_clk),
    .D(_0735_),
    .RESET_B(_0206_),
    .Q(\output_c[4][21] ));
 sky130_fd_sc_hd__dfrtp_1 _4971_ (.CLK(clknet_leaf_32_clk),
    .D(_0736_),
    .RESET_B(_0207_),
    .Q(\output_c[4][22] ));
 sky130_fd_sc_hd__dfrtp_1 _4972_ (.CLK(clknet_leaf_32_clk),
    .D(_0737_),
    .RESET_B(_0208_),
    .Q(\output_c[4][23] ));
 sky130_fd_sc_hd__dfrtp_1 _4973_ (.CLK(clknet_leaf_32_clk),
    .D(_0738_),
    .RESET_B(_0209_),
    .Q(\output_c[4][24] ));
 sky130_fd_sc_hd__dfrtp_1 _4974_ (.CLK(clknet_leaf_32_clk),
    .D(_0739_),
    .RESET_B(_0210_),
    .Q(\output_c[4][25] ));
 sky130_fd_sc_hd__dfrtp_1 _4975_ (.CLK(clknet_leaf_33_clk),
    .D(_0740_),
    .RESET_B(_0211_),
    .Q(\output_c[4][26] ));
 sky130_fd_sc_hd__dfrtp_1 _4976_ (.CLK(clknet_leaf_32_clk),
    .D(_0741_),
    .RESET_B(_0212_),
    .Q(\output_c[4][27] ));
 sky130_fd_sc_hd__dfrtp_1 _4977_ (.CLK(clknet_leaf_32_clk),
    .D(_0742_),
    .RESET_B(_0213_),
    .Q(\output_c[4][28] ));
 sky130_fd_sc_hd__dfrtp_1 _4978_ (.CLK(clknet_leaf_32_clk),
    .D(_0743_),
    .RESET_B(_0214_),
    .Q(\output_c[4][29] ));
 sky130_fd_sc_hd__dfrtp_1 _4979_ (.CLK(clknet_leaf_34_clk),
    .D(_0744_),
    .RESET_B(_0215_),
    .Q(\output_c[4][30] ));
 sky130_fd_sc_hd__dfrtp_1 _4980_ (.CLK(clknet_leaf_34_clk),
    .D(_0745_),
    .RESET_B(_0216_),
    .Q(\output_c[4][31] ));
 sky130_fd_sc_hd__dfrtp_1 _4981_ (.CLK(clknet_leaf_36_clk),
    .D(_0746_),
    .RESET_B(_0217_),
    .Q(\output_c[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _4982_ (.CLK(clknet_leaf_36_clk),
    .D(_0747_),
    .RESET_B(_0218_),
    .Q(\output_c[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _4983_ (.CLK(clknet_leaf_36_clk),
    .D(_0748_),
    .RESET_B(_0219_),
    .Q(\output_c[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _4984_ (.CLK(clknet_leaf_34_clk),
    .D(_0749_),
    .RESET_B(_0220_),
    .Q(\output_c[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _4985_ (.CLK(clknet_leaf_34_clk),
    .D(_0750_),
    .RESET_B(_0221_),
    .Q(\output_c[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _4986_ (.CLK(clknet_leaf_34_clk),
    .D(_0751_),
    .RESET_B(_0222_),
    .Q(\output_c[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _4987_ (.CLK(clknet_leaf_32_clk),
    .D(_0752_),
    .RESET_B(_0223_),
    .Q(\output_c[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _4988_ (.CLK(clknet_leaf_34_clk),
    .D(_0753_),
    .RESET_B(_0224_),
    .Q(\output_c[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _4989_ (.CLK(clknet_leaf_33_clk),
    .D(_0754_),
    .RESET_B(_0225_),
    .Q(\output_c[5][8] ));
 sky130_fd_sc_hd__dfrtp_1 _4990_ (.CLK(clknet_leaf_33_clk),
    .D(_0755_),
    .RESET_B(_0226_),
    .Q(\output_c[5][9] ));
 sky130_fd_sc_hd__dfrtp_1 _4991_ (.CLK(clknet_leaf_33_clk),
    .D(_0756_),
    .RESET_B(_0227_),
    .Q(\output_c[5][10] ));
 sky130_fd_sc_hd__dfrtp_1 _4992_ (.CLK(clknet_leaf_33_clk),
    .D(_0757_),
    .RESET_B(_0228_),
    .Q(\output_c[5][11] ));
 sky130_fd_sc_hd__dfrtp_1 _4993_ (.CLK(clknet_leaf_32_clk),
    .D(_0758_),
    .RESET_B(_0229_),
    .Q(\output_c[5][12] ));
 sky130_fd_sc_hd__dfrtp_1 _4994_ (.CLK(clknet_leaf_33_clk),
    .D(_0759_),
    .RESET_B(_0230_),
    .Q(\output_c[5][13] ));
 sky130_fd_sc_hd__dfrtp_1 _4995_ (.CLK(clknet_leaf_33_clk),
    .D(_0760_),
    .RESET_B(_0231_),
    .Q(\output_c[5][14] ));
 sky130_fd_sc_hd__dfrtp_1 _4996_ (.CLK(clknet_leaf_33_clk),
    .D(_0761_),
    .RESET_B(_0232_),
    .Q(\output_c[5][15] ));
 sky130_fd_sc_hd__dfrtp_1 _4997_ (.CLK(clknet_leaf_38_clk),
    .D(_0762_),
    .RESET_B(_0233_),
    .Q(\output_c[5][16] ));
 sky130_fd_sc_hd__dfrtp_1 _4998_ (.CLK(clknet_leaf_38_clk),
    .D(_0763_),
    .RESET_B(_0234_),
    .Q(\output_c[5][17] ));
 sky130_fd_sc_hd__dfrtp_1 _4999_ (.CLK(clknet_leaf_38_clk),
    .D(_0764_),
    .RESET_B(_0235_),
    .Q(\output_c[5][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5000_ (.CLK(clknet_leaf_38_clk),
    .D(_0765_),
    .RESET_B(_0236_),
    .Q(\output_c[5][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5001_ (.CLK(clknet_leaf_38_clk),
    .D(_0766_),
    .RESET_B(_0237_),
    .Q(\output_c[5][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5002_ (.CLK(clknet_leaf_38_clk),
    .D(_0767_),
    .RESET_B(_0238_),
    .Q(\output_c[5][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5003_ (.CLK(clknet_leaf_38_clk),
    .D(_0768_),
    .RESET_B(_0239_),
    .Q(\output_c[5][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5004_ (.CLK(clknet_leaf_38_clk),
    .D(_0769_),
    .RESET_B(_0240_),
    .Q(\output_c[5][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5005_ (.CLK(clknet_leaf_38_clk),
    .D(_0770_),
    .RESET_B(_0241_),
    .Q(\output_c[5][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5006_ (.CLK(clknet_leaf_37_clk),
    .D(_0771_),
    .RESET_B(_0242_),
    .Q(\output_c[5][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5007_ (.CLK(clknet_leaf_37_clk),
    .D(_0772_),
    .RESET_B(_0243_),
    .Q(\output_c[5][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5008_ (.CLK(clknet_leaf_34_clk),
    .D(_0773_),
    .RESET_B(_0244_),
    .Q(\output_c[5][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5009_ (.CLK(clknet_leaf_34_clk),
    .D(_0774_),
    .RESET_B(_0245_),
    .Q(\output_c[5][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5010_ (.CLK(clknet_leaf_37_clk),
    .D(net317),
    .RESET_B(_0246_),
    .Q(\output_c[5][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5011_ (.CLK(clknet_leaf_37_clk),
    .D(_0776_),
    .RESET_B(_0247_),
    .Q(\output_c[5][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5012_ (.CLK(clknet_leaf_37_clk),
    .D(_0777_),
    .RESET_B(_0248_),
    .Q(\output_c[5][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5013_ (.CLK(clknet_leaf_36_clk),
    .D(_0778_),
    .RESET_B(_0249_),
    .Q(\output_c[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5014_ (.CLK(clknet_leaf_37_clk),
    .D(_0779_),
    .RESET_B(_0250_),
    .Q(\output_c[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5015_ (.CLK(clknet_leaf_37_clk),
    .D(net451),
    .RESET_B(_0251_),
    .Q(\output_c[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5016_ (.CLK(clknet_leaf_37_clk),
    .D(_0781_),
    .RESET_B(_0252_),
    .Q(\output_c[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5017_ (.CLK(clknet_leaf_0_clk),
    .D(_0782_),
    .RESET_B(_0253_),
    .Q(\output_c[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5018_ (.CLK(clknet_leaf_0_clk),
    .D(_0783_),
    .RESET_B(_0254_),
    .Q(\output_c[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5019_ (.CLK(clknet_leaf_39_clk),
    .D(_0784_),
    .RESET_B(_0255_),
    .Q(\output_c[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5020_ (.CLK(clknet_leaf_40_clk),
    .D(_0785_),
    .RESET_B(_0256_),
    .Q(\output_c[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5021_ (.CLK(clknet_leaf_40_clk),
    .D(_0786_),
    .RESET_B(_0257_),
    .Q(\output_c[6][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5022_ (.CLK(clknet_leaf_40_clk),
    .D(_0787_),
    .RESET_B(_0258_),
    .Q(\output_c[6][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5023_ (.CLK(clknet_leaf_40_clk),
    .D(_0788_),
    .RESET_B(_0259_),
    .Q(\output_c[6][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5024_ (.CLK(clknet_leaf_40_clk),
    .D(_0789_),
    .RESET_B(_0260_),
    .Q(\output_c[6][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5025_ (.CLK(clknet_leaf_40_clk),
    .D(_0790_),
    .RESET_B(_0261_),
    .Q(\output_c[6][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5026_ (.CLK(clknet_leaf_0_clk),
    .D(_0791_),
    .RESET_B(_0262_),
    .Q(\output_c[6][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5027_ (.CLK(clknet_leaf_41_clk),
    .D(_0792_),
    .RESET_B(_0263_),
    .Q(\output_c[6][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5028_ (.CLK(clknet_leaf_41_clk),
    .D(_0793_),
    .RESET_B(_0264_),
    .Q(\output_c[6][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5029_ (.CLK(clknet_leaf_41_clk),
    .D(_0794_),
    .RESET_B(_0265_),
    .Q(\output_c[6][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5030_ (.CLK(clknet_leaf_40_clk),
    .D(_0795_),
    .RESET_B(_0266_),
    .Q(\output_c[6][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5031_ (.CLK(clknet_leaf_41_clk),
    .D(_0796_),
    .RESET_B(_0267_),
    .Q(\output_c[6][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5032_ (.CLK(clknet_leaf_41_clk),
    .D(_0797_),
    .RESET_B(_0268_),
    .Q(\output_c[6][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5033_ (.CLK(clknet_leaf_41_clk),
    .D(_0798_),
    .RESET_B(_0269_),
    .Q(\output_c[6][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5034_ (.CLK(clknet_leaf_41_clk),
    .D(_0799_),
    .RESET_B(_0270_),
    .Q(\output_c[6][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5035_ (.CLK(clknet_leaf_41_clk),
    .D(_0800_),
    .RESET_B(_0271_),
    .Q(\output_c[6][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5036_ (.CLK(clknet_leaf_41_clk),
    .D(_0801_),
    .RESET_B(_0272_),
    .Q(\output_c[6][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5037_ (.CLK(clknet_leaf_0_clk),
    .D(_0802_),
    .RESET_B(_0273_),
    .Q(\output_c[6][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5038_ (.CLK(clknet_leaf_0_clk),
    .D(_0803_),
    .RESET_B(_0274_),
    .Q(\output_c[6][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5039_ (.CLK(clknet_leaf_0_clk),
    .D(_0804_),
    .RESET_B(_0275_),
    .Q(\output_c[6][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5040_ (.CLK(clknet_leaf_0_clk),
    .D(_0805_),
    .RESET_B(_0276_),
    .Q(\output_c[6][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5041_ (.CLK(clknet_leaf_0_clk),
    .D(_0806_),
    .RESET_B(_0277_),
    .Q(\output_c[6][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5042_ (.CLK(clknet_leaf_0_clk),
    .D(_0807_),
    .RESET_B(_0278_),
    .Q(\output_c[6][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5043_ (.CLK(clknet_leaf_0_clk),
    .D(_0808_),
    .RESET_B(_0279_),
    .Q(\output_c[6][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5044_ (.CLK(clknet_leaf_3_clk),
    .D(_0809_),
    .RESET_B(_0280_),
    .Q(\output_c[6][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5045_ (.CLK(clknet_leaf_4_clk),
    .D(_0810_),
    .RESET_B(_0281_),
    .Q(\output_c[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5046_ (.CLK(clknet_leaf_37_clk),
    .D(_0811_),
    .RESET_B(_0282_),
    .Q(\output_c[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5047_ (.CLK(clknet_leaf_37_clk),
    .D(_0812_),
    .RESET_B(_0283_),
    .Q(\output_c[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5048_ (.CLK(clknet_leaf_37_clk),
    .D(_0813_),
    .RESET_B(_0284_),
    .Q(\output_c[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5049_ (.CLK(clknet_leaf_37_clk),
    .D(_0814_),
    .RESET_B(_0285_),
    .Q(\output_c[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5050_ (.CLK(clknet_leaf_39_clk),
    .D(_0815_),
    .RESET_B(_0286_),
    .Q(\output_c[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5051_ (.CLK(clknet_leaf_39_clk),
    .D(_0816_),
    .RESET_B(_0287_),
    .Q(\output_c[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5052_ (.CLK(clknet_leaf_39_clk),
    .D(_0817_),
    .RESET_B(_0288_),
    .Q(\output_c[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5053_ (.CLK(clknet_leaf_39_clk),
    .D(_0818_),
    .RESET_B(_0289_),
    .Q(\output_c[7][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5054_ (.CLK(clknet_leaf_39_clk),
    .D(_0819_),
    .RESET_B(_0290_),
    .Q(\output_c[7][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5055_ (.CLK(clknet_leaf_39_clk),
    .D(_0820_),
    .RESET_B(_0291_),
    .Q(\output_c[7][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5056_ (.CLK(clknet_leaf_40_clk),
    .D(_0821_),
    .RESET_B(_0292_),
    .Q(\output_c[7][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5057_ (.CLK(clknet_leaf_40_clk),
    .D(_0822_),
    .RESET_B(_0293_),
    .Q(\output_c[7][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5058_ (.CLK(clknet_leaf_40_clk),
    .D(_0823_),
    .RESET_B(_0294_),
    .Q(\output_c[7][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5059_ (.CLK(clknet_leaf_40_clk),
    .D(_0824_),
    .RESET_B(_0295_),
    .Q(\output_c[7][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5060_ (.CLK(clknet_leaf_39_clk),
    .D(_0825_),
    .RESET_B(_0296_),
    .Q(\output_c[7][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5061_ (.CLK(clknet_leaf_39_clk),
    .D(_0826_),
    .RESET_B(_0297_),
    .Q(\output_c[7][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5062_ (.CLK(clknet_leaf_39_clk),
    .D(_0827_),
    .RESET_B(_0298_),
    .Q(\output_c[7][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5063_ (.CLK(clknet_leaf_39_clk),
    .D(_0828_),
    .RESET_B(_0299_),
    .Q(\output_c[7][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5064_ (.CLK(clknet_leaf_38_clk),
    .D(_0829_),
    .RESET_B(_0300_),
    .Q(\output_c[7][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5065_ (.CLK(clknet_leaf_38_clk),
    .D(_0830_),
    .RESET_B(_0301_),
    .Q(\output_c[7][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5066_ (.CLK(clknet_leaf_38_clk),
    .D(_0831_),
    .RESET_B(_0302_),
    .Q(\output_c[7][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5067_ (.CLK(clknet_leaf_38_clk),
    .D(_0832_),
    .RESET_B(_0303_),
    .Q(\output_c[7][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5068_ (.CLK(clknet_leaf_38_clk),
    .D(_0833_),
    .RESET_B(_0304_),
    .Q(\output_c[7][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5069_ (.CLK(clknet_leaf_39_clk),
    .D(_0834_),
    .RESET_B(_0305_),
    .Q(\output_c[7][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5070_ (.CLK(clknet_leaf_39_clk),
    .D(_0835_),
    .RESET_B(_0306_),
    .Q(\output_c[7][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5071_ (.CLK(clknet_leaf_38_clk),
    .D(_0836_),
    .RESET_B(_0307_),
    .Q(\output_c[7][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5072_ (.CLK(clknet_leaf_37_clk),
    .D(_0837_),
    .RESET_B(_0308_),
    .Q(\output_c[7][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5073_ (.CLK(clknet_leaf_37_clk),
    .D(_0838_),
    .RESET_B(_0309_),
    .Q(\output_c[7][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5074_ (.CLK(clknet_leaf_37_clk),
    .D(_0839_),
    .RESET_B(_0310_),
    .Q(\output_c[7][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5075_ (.CLK(clknet_leaf_37_clk),
    .D(_0840_),
    .RESET_B(_0311_),
    .Q(\output_c[7][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5076_ (.CLK(clknet_leaf_37_clk),
    .D(_0841_),
    .RESET_B(_0312_),
    .Q(\output_c[7][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5077_ (.CLK(clknet_leaf_36_clk),
    .D(_0842_),
    .RESET_B(_0313_),
    .Q(\output_c[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5078_ (.CLK(clknet_leaf_36_clk),
    .D(_0843_),
    .RESET_B(_0314_),
    .Q(\output_c[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5079_ (.CLK(clknet_leaf_36_clk),
    .D(net429),
    .RESET_B(_0315_),
    .Q(\output_c[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5080_ (.CLK(clknet_leaf_36_clk),
    .D(_0845_),
    .RESET_B(_0316_),
    .Q(\output_c[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5081_ (.CLK(clknet_leaf_36_clk),
    .D(_0846_),
    .RESET_B(_0317_),
    .Q(\output_c[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5082_ (.CLK(clknet_leaf_36_clk),
    .D(_0847_),
    .RESET_B(_0318_),
    .Q(\output_c[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5083_ (.CLK(clknet_leaf_35_clk),
    .D(_0848_),
    .RESET_B(_0319_),
    .Q(\output_c[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5084_ (.CLK(clknet_leaf_35_clk),
    .D(_0849_),
    .RESET_B(_0320_),
    .Q(\output_c[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5085_ (.CLK(clknet_leaf_35_clk),
    .D(_0850_),
    .RESET_B(_0321_),
    .Q(\output_c[8][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5086_ (.CLK(clknet_leaf_34_clk),
    .D(_0851_),
    .RESET_B(_0322_),
    .Q(\output_c[8][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5087_ (.CLK(clknet_leaf_34_clk),
    .D(_0852_),
    .RESET_B(_0323_),
    .Q(\output_c[8][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5088_ (.CLK(clknet_leaf_34_clk),
    .D(_0853_),
    .RESET_B(_0324_),
    .Q(\output_c[8][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5089_ (.CLK(clknet_leaf_34_clk),
    .D(_0854_),
    .RESET_B(_0325_),
    .Q(\output_c[8][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5090_ (.CLK(clknet_leaf_32_clk),
    .D(_0855_),
    .RESET_B(_0326_),
    .Q(\output_c[8][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5091_ (.CLK(clknet_leaf_34_clk),
    .D(_0856_),
    .RESET_B(_0327_),
    .Q(\output_c[8][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5092_ (.CLK(clknet_leaf_35_clk),
    .D(_0857_),
    .RESET_B(_0328_),
    .Q(\output_c[8][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5093_ (.CLK(clknet_leaf_35_clk),
    .D(_0858_),
    .RESET_B(_0329_),
    .Q(\output_c[8][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5094_ (.CLK(clknet_leaf_35_clk),
    .D(_0859_),
    .RESET_B(_0330_),
    .Q(\output_c[8][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5095_ (.CLK(clknet_leaf_35_clk),
    .D(_0860_),
    .RESET_B(_0331_),
    .Q(\output_c[8][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5096_ (.CLK(clknet_leaf_27_clk),
    .D(_0861_),
    .RESET_B(_0332_),
    .Q(\output_c[8][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5097_ (.CLK(clknet_leaf_27_clk),
    .D(_0862_),
    .RESET_B(_0333_),
    .Q(\output_c[8][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5098_ (.CLK(clknet_leaf_27_clk),
    .D(_0863_),
    .RESET_B(_0334_),
    .Q(\output_c[8][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5099_ (.CLK(clknet_leaf_27_clk),
    .D(_0864_),
    .RESET_B(_0335_),
    .Q(\output_c[8][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5100_ (.CLK(clknet_leaf_35_clk),
    .D(_0865_),
    .RESET_B(_0336_),
    .Q(\output_c[8][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5101_ (.CLK(clknet_leaf_36_clk),
    .D(_0866_),
    .RESET_B(_0337_),
    .Q(\output_c[8][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5102_ (.CLK(clknet_leaf_36_clk),
    .D(_0867_),
    .RESET_B(_0338_),
    .Q(\output_c[8][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5103_ (.CLK(clknet_leaf_27_clk),
    .D(_0868_),
    .RESET_B(_0339_),
    .Q(\output_c[8][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5104_ (.CLK(clknet_leaf_27_clk),
    .D(_0869_),
    .RESET_B(_0340_),
    .Q(\output_c[8][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5105_ (.CLK(clknet_leaf_26_clk),
    .D(_0870_),
    .RESET_B(_0341_),
    .Q(\output_c[8][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5106_ (.CLK(clknet_leaf_26_clk),
    .D(_0871_),
    .RESET_B(_0342_),
    .Q(\output_c[8][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5107_ (.CLK(clknet_leaf_26_clk),
    .D(_0872_),
    .RESET_B(_0343_),
    .Q(\output_c[8][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5108_ (.CLK(clknet_leaf_26_clk),
    .D(_0873_),
    .RESET_B(_0344_),
    .Q(\output_c[8][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5109_ (.CLK(clknet_leaf_26_clk),
    .D(_0874_),
    .RESET_B(_0345_),
    .Q(\output_c[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5110_ (.CLK(clknet_leaf_26_clk),
    .D(_0875_),
    .RESET_B(_0346_),
    .Q(\output_c[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5111_ (.CLK(clknet_leaf_25_clk),
    .D(net447),
    .RESET_B(_0347_),
    .Q(\output_c[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5112_ (.CLK(clknet_leaf_26_clk),
    .D(net198),
    .RESET_B(_0348_),
    .Q(\output_c[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5113_ (.CLK(clknet_leaf_24_clk),
    .D(_0878_),
    .RESET_B(_0349_),
    .Q(\output_c[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5114_ (.CLK(clknet_leaf_24_clk),
    .D(_0879_),
    .RESET_B(_0350_),
    .Q(\output_c[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5115_ (.CLK(clknet_leaf_24_clk),
    .D(_0880_),
    .RESET_B(_0351_),
    .Q(\output_c[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5116_ (.CLK(clknet_leaf_23_clk),
    .D(_0881_),
    .RESET_B(_0352_),
    .Q(\output_c[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5117_ (.CLK(clknet_leaf_23_clk),
    .D(_0882_),
    .RESET_B(_0353_),
    .Q(\output_c[9][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5118_ (.CLK(clknet_leaf_23_clk),
    .D(_0883_),
    .RESET_B(_0354_),
    .Q(\output_c[9][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5119_ (.CLK(clknet_leaf_23_clk),
    .D(_0884_),
    .RESET_B(_0355_),
    .Q(\output_c[9][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5120_ (.CLK(clknet_leaf_23_clk),
    .D(_0885_),
    .RESET_B(_0356_),
    .Q(\output_c[9][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5121_ (.CLK(clknet_leaf_22_clk),
    .D(_0886_),
    .RESET_B(_0357_),
    .Q(\output_c[9][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5122_ (.CLK(clknet_leaf_22_clk),
    .D(_0887_),
    .RESET_B(_0358_),
    .Q(\output_c[9][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5123_ (.CLK(clknet_leaf_22_clk),
    .D(_0888_),
    .RESET_B(_0359_),
    .Q(\output_c[9][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5124_ (.CLK(clknet_leaf_22_clk),
    .D(_0889_),
    .RESET_B(_0360_),
    .Q(\output_c[9][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5125_ (.CLK(clknet_leaf_21_clk),
    .D(_0890_),
    .RESET_B(_0361_),
    .Q(\output_c[9][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5126_ (.CLK(clknet_leaf_22_clk),
    .D(_0891_),
    .RESET_B(_0362_),
    .Q(\output_c[9][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5127_ (.CLK(clknet_leaf_22_clk),
    .D(_0892_),
    .RESET_B(_0363_),
    .Q(\output_c[9][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5128_ (.CLK(clknet_leaf_21_clk),
    .D(_0893_),
    .RESET_B(_0364_),
    .Q(\output_c[9][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5129_ (.CLK(clknet_leaf_21_clk),
    .D(_0894_),
    .RESET_B(_0365_),
    .Q(\output_c[9][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5130_ (.CLK(clknet_leaf_21_clk),
    .D(_0895_),
    .RESET_B(_0366_),
    .Q(\output_c[9][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5131_ (.CLK(clknet_leaf_21_clk),
    .D(_0896_),
    .RESET_B(_0367_),
    .Q(\output_c[9][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5132_ (.CLK(clknet_leaf_21_clk),
    .D(_0897_),
    .RESET_B(_0368_),
    .Q(\output_c[9][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5133_ (.CLK(clknet_leaf_20_clk),
    .D(_0898_),
    .RESET_B(_0369_),
    .Q(\output_c[9][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5134_ (.CLK(clknet_leaf_19_clk),
    .D(_0899_),
    .RESET_B(_0370_),
    .Q(\output_c[9][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5135_ (.CLK(clknet_leaf_20_clk),
    .D(_0900_),
    .RESET_B(_0371_),
    .Q(\output_c[9][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5136_ (.CLK(clknet_leaf_19_clk),
    .D(_0901_),
    .RESET_B(_0372_),
    .Q(\output_c[9][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5137_ (.CLK(clknet_leaf_21_clk),
    .D(_0902_),
    .RESET_B(_0373_),
    .Q(\output_c[9][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5138_ (.CLK(clknet_leaf_19_clk),
    .D(net319),
    .RESET_B(_0374_),
    .Q(\output_c[9][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5139_ (.CLK(clknet_leaf_19_clk),
    .D(_0904_),
    .RESET_B(_0375_),
    .Q(\output_c[9][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5140_ (.CLK(clknet_leaf_19_clk),
    .D(_0905_),
    .RESET_B(_0376_),
    .Q(\output_c[9][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5141_ (.CLK(clknet_leaf_15_clk),
    .D(_0906_),
    .RESET_B(_0377_),
    .Q(\output_c[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5142_ (.CLK(clknet_leaf_16_clk),
    .D(_0907_),
    .RESET_B(_0378_),
    .Q(\output_c[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5143_ (.CLK(clknet_leaf_16_clk),
    .D(_0908_),
    .RESET_B(_0379_),
    .Q(\output_c[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5144_ (.CLK(clknet_leaf_16_clk),
    .D(_0909_),
    .RESET_B(_0380_),
    .Q(\output_c[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5145_ (.CLK(clknet_leaf_16_clk),
    .D(_0910_),
    .RESET_B(_0381_),
    .Q(\output_c[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5146_ (.CLK(clknet_leaf_16_clk),
    .D(_0911_),
    .RESET_B(_0382_),
    .Q(\output_c[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5147_ (.CLK(clknet_leaf_19_clk),
    .D(_0912_),
    .RESET_B(_0383_),
    .Q(\output_c[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5148_ (.CLK(clknet_leaf_19_clk),
    .D(_0913_),
    .RESET_B(_0384_),
    .Q(\output_c[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5149_ (.CLK(clknet_leaf_18_clk),
    .D(_0914_),
    .RESET_B(_0385_),
    .Q(\output_c[10][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5150_ (.CLK(clknet_leaf_18_clk),
    .D(_0915_),
    .RESET_B(_0386_),
    .Q(\output_c[10][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5151_ (.CLK(clknet_leaf_19_clk),
    .D(_0916_),
    .RESET_B(_0387_),
    .Q(\output_c[10][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5152_ (.CLK(clknet_leaf_19_clk),
    .D(_0917_),
    .RESET_B(_0388_),
    .Q(\output_c[10][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5153_ (.CLK(clknet_leaf_20_clk),
    .D(_0918_),
    .RESET_B(_0389_),
    .Q(\output_c[10][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5154_ (.CLK(clknet_leaf_19_clk),
    .D(_0919_),
    .RESET_B(_0390_),
    .Q(\output_c[10][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5155_ (.CLK(clknet_leaf_20_clk),
    .D(_0920_),
    .RESET_B(_0391_),
    .Q(\output_c[10][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5156_ (.CLK(clknet_leaf_20_clk),
    .D(_0921_),
    .RESET_B(_0392_),
    .Q(\output_c[10][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5157_ (.CLK(clknet_leaf_18_clk),
    .D(_0922_),
    .RESET_B(_0393_),
    .Q(\output_c[10][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5158_ (.CLK(clknet_leaf_19_clk),
    .D(_0923_),
    .RESET_B(_0394_),
    .Q(\output_c[10][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5159_ (.CLK(clknet_leaf_18_clk),
    .D(_0924_),
    .RESET_B(_0395_),
    .Q(\output_c[10][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5160_ (.CLK(clknet_leaf_18_clk),
    .D(_0925_),
    .RESET_B(_0396_),
    .Q(\output_c[10][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5161_ (.CLK(clknet_leaf_18_clk),
    .D(_0926_),
    .RESET_B(_0397_),
    .Q(\output_c[10][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5162_ (.CLK(clknet_leaf_18_clk),
    .D(_0927_),
    .RESET_B(_0398_),
    .Q(\output_c[10][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5163_ (.CLK(clknet_leaf_18_clk),
    .D(_0928_),
    .RESET_B(_0399_),
    .Q(\output_c[10][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5164_ (.CLK(clknet_leaf_18_clk),
    .D(_0929_),
    .RESET_B(_0400_),
    .Q(\output_c[10][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5165_ (.CLK(clknet_leaf_18_clk),
    .D(_0930_),
    .RESET_B(_0401_),
    .Q(\output_c[10][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5166_ (.CLK(clknet_leaf_17_clk),
    .D(_0931_),
    .RESET_B(_0402_),
    .Q(\output_c[10][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5167_ (.CLK(clknet_leaf_17_clk),
    .D(_0932_),
    .RESET_B(_0403_),
    .Q(\output_c[10][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5168_ (.CLK(clknet_leaf_17_clk),
    .D(_0933_),
    .RESET_B(_0404_),
    .Q(\output_c[10][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5169_ (.CLK(clknet_leaf_17_clk),
    .D(_0934_),
    .RESET_B(_0405_),
    .Q(\output_c[10][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5170_ (.CLK(clknet_leaf_17_clk),
    .D(_0935_),
    .RESET_B(_0406_),
    .Q(\output_c[10][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5171_ (.CLK(clknet_leaf_17_clk),
    .D(_0936_),
    .RESET_B(_0407_),
    .Q(\output_c[10][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5172_ (.CLK(clknet_leaf_12_clk),
    .D(_0937_),
    .RESET_B(_0408_),
    .Q(\output_c[10][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5173_ (.CLK(clknet_leaf_14_clk),
    .D(_0938_),
    .RESET_B(_0409_),
    .Q(\output_c[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5174_ (.CLK(clknet_leaf_14_clk),
    .D(_0939_),
    .RESET_B(_0410_),
    .Q(\output_c[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5175_ (.CLK(clknet_leaf_14_clk),
    .D(net425),
    .RESET_B(_0411_),
    .Q(\output_c[11][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5176_ (.CLK(clknet_leaf_14_clk),
    .D(_0941_),
    .RESET_B(_0412_),
    .Q(\output_c[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5177_ (.CLK(clknet_leaf_13_clk),
    .D(_0942_),
    .RESET_B(_0413_),
    .Q(\output_c[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5178_ (.CLK(clknet_leaf_13_clk),
    .D(_0943_),
    .RESET_B(_0414_),
    .Q(\output_c[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5179_ (.CLK(clknet_leaf_12_clk),
    .D(_0944_),
    .RESET_B(_0415_),
    .Q(\output_c[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5180_ (.CLK(clknet_leaf_12_clk),
    .D(_0945_),
    .RESET_B(_0416_),
    .Q(\output_c[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5181_ (.CLK(clknet_leaf_12_clk),
    .D(_0946_),
    .RESET_B(_0417_),
    .Q(\output_c[11][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5182_ (.CLK(clknet_leaf_12_clk),
    .D(_0947_),
    .RESET_B(_0418_),
    .Q(\output_c[11][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5183_ (.CLK(clknet_leaf_12_clk),
    .D(_0948_),
    .RESET_B(_0419_),
    .Q(\output_c[11][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5184_ (.CLK(clknet_leaf_12_clk),
    .D(_0949_),
    .RESET_B(_0420_),
    .Q(\output_c[11][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5185_ (.CLK(clknet_leaf_12_clk),
    .D(_0950_),
    .RESET_B(_0421_),
    .Q(\output_c[11][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5186_ (.CLK(clknet_leaf_12_clk),
    .D(_0951_),
    .RESET_B(_0422_),
    .Q(\output_c[11][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5187_ (.CLK(clknet_leaf_12_clk),
    .D(_0952_),
    .RESET_B(_0423_),
    .Q(\output_c[11][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5188_ (.CLK(clknet_leaf_12_clk),
    .D(_0953_),
    .RESET_B(_0424_),
    .Q(\output_c[11][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5189_ (.CLK(clknet_leaf_12_clk),
    .D(_0954_),
    .RESET_B(_0425_),
    .Q(\output_c[11][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5190_ (.CLK(clknet_leaf_11_clk),
    .D(_0955_),
    .RESET_B(_0426_),
    .Q(\output_c[11][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5191_ (.CLK(clknet_leaf_11_clk),
    .D(_0956_),
    .RESET_B(_0427_),
    .Q(\output_c[11][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5192_ (.CLK(clknet_leaf_10_clk),
    .D(_0957_),
    .RESET_B(_0428_),
    .Q(\output_c[11][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5193_ (.CLK(clknet_leaf_10_clk),
    .D(_0958_),
    .RESET_B(_0429_),
    .Q(\output_c[11][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5194_ (.CLK(clknet_leaf_10_clk),
    .D(_0959_),
    .RESET_B(_0430_),
    .Q(\output_c[11][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5195_ (.CLK(clknet_leaf_10_clk),
    .D(_0960_),
    .RESET_B(_0431_),
    .Q(\output_c[11][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5196_ (.CLK(clknet_leaf_11_clk),
    .D(_0961_),
    .RESET_B(_0432_),
    .Q(\output_c[11][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5197_ (.CLK(clknet_leaf_11_clk),
    .D(_0962_),
    .RESET_B(_0433_),
    .Q(\output_c[11][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5198_ (.CLK(clknet_leaf_11_clk),
    .D(_0963_),
    .RESET_B(_0434_),
    .Q(\output_c[11][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5199_ (.CLK(clknet_leaf_11_clk),
    .D(_0964_),
    .RESET_B(_0435_),
    .Q(\output_c[11][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5200_ (.CLK(clknet_leaf_11_clk),
    .D(_0965_),
    .RESET_B(_0436_),
    .Q(\output_c[11][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5201_ (.CLK(clknet_leaf_14_clk),
    .D(_0966_),
    .RESET_B(_0437_),
    .Q(\output_c[11][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5202_ (.CLK(clknet_leaf_14_clk),
    .D(_0967_),
    .RESET_B(_0438_),
    .Q(\output_c[11][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5203_ (.CLK(clknet_leaf_13_clk),
    .D(_0968_),
    .RESET_B(_0439_),
    .Q(\output_c[11][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5204_ (.CLK(clknet_leaf_14_clk),
    .D(_0969_),
    .RESET_B(_0440_),
    .Q(\output_c[11][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5205_ (.CLK(clknet_leaf_14_clk),
    .D(_0970_),
    .RESET_B(_0441_),
    .Q(\output_c[12][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5206_ (.CLK(clknet_leaf_14_clk),
    .D(_0971_),
    .RESET_B(_0442_),
    .Q(\output_c[12][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5207_ (.CLK(clknet_leaf_14_clk),
    .D(_0972_),
    .RESET_B(_0443_),
    .Q(\output_c[12][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5208_ (.CLK(clknet_leaf_14_clk),
    .D(_0973_),
    .RESET_B(_0444_),
    .Q(\output_c[12][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5209_ (.CLK(clknet_leaf_5_clk),
    .D(_0974_),
    .RESET_B(_0445_),
    .Q(\output_c[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5210_ (.CLK(clknet_leaf_11_clk),
    .D(_0975_),
    .RESET_B(_0446_),
    .Q(\output_c[12][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5211_ (.CLK(clknet_leaf_11_clk),
    .D(_0976_),
    .RESET_B(_0447_),
    .Q(\output_c[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5212_ (.CLK(clknet_leaf_10_clk),
    .D(_0977_),
    .RESET_B(_0448_),
    .Q(\output_c[12][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5213_ (.CLK(clknet_leaf_8_clk),
    .D(_0978_),
    .RESET_B(_0449_),
    .Q(\output_c[12][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5214_ (.CLK(clknet_leaf_10_clk),
    .D(_0979_),
    .RESET_B(_0450_),
    .Q(\output_c[12][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5215_ (.CLK(clknet_leaf_10_clk),
    .D(_0980_),
    .RESET_B(_0451_),
    .Q(\output_c[12][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5216_ (.CLK(clknet_leaf_10_clk),
    .D(_0981_),
    .RESET_B(_0452_),
    .Q(\output_c[12][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5217_ (.CLK(clknet_leaf_10_clk),
    .D(_0982_),
    .RESET_B(_0453_),
    .Q(\output_c[12][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5218_ (.CLK(clknet_leaf_9_clk),
    .D(_0983_),
    .RESET_B(_0454_),
    .Q(\output_c[12][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5219_ (.CLK(clknet_leaf_10_clk),
    .D(_0984_),
    .RESET_B(_0455_),
    .Q(\output_c[12][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5220_ (.CLK(clknet_leaf_9_clk),
    .D(_0985_),
    .RESET_B(_0456_),
    .Q(\output_c[12][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5221_ (.CLK(clknet_leaf_9_clk),
    .D(_0986_),
    .RESET_B(_0457_),
    .Q(\output_c[12][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5222_ (.CLK(clknet_leaf_9_clk),
    .D(_0987_),
    .RESET_B(_0458_),
    .Q(\output_c[12][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5223_ (.CLK(clknet_leaf_9_clk),
    .D(_0988_),
    .RESET_B(_0459_),
    .Q(\output_c[12][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5224_ (.CLK(clknet_leaf_9_clk),
    .D(_0989_),
    .RESET_B(_0460_),
    .Q(\output_c[12][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5225_ (.CLK(clknet_leaf_9_clk),
    .D(_0990_),
    .RESET_B(_0461_),
    .Q(\output_c[12][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5226_ (.CLK(clknet_leaf_8_clk),
    .D(_0991_),
    .RESET_B(_0462_),
    .Q(\output_c[12][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5227_ (.CLK(clknet_leaf_8_clk),
    .D(_0992_),
    .RESET_B(_0463_),
    .Q(\output_c[12][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5228_ (.CLK(clknet_leaf_8_clk),
    .D(_0993_),
    .RESET_B(_0464_),
    .Q(\output_c[12][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5229_ (.CLK(clknet_leaf_8_clk),
    .D(_0994_),
    .RESET_B(_0465_),
    .Q(\output_c[12][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5230_ (.CLK(clknet_leaf_8_clk),
    .D(_0995_),
    .RESET_B(_0466_),
    .Q(\output_c[12][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5231_ (.CLK(clknet_leaf_8_clk),
    .D(_0996_),
    .RESET_B(_0467_),
    .Q(\output_c[12][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5232_ (.CLK(clknet_leaf_8_clk),
    .D(_0997_),
    .RESET_B(_0468_),
    .Q(\output_c[12][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5233_ (.CLK(clknet_leaf_10_clk),
    .D(_0998_),
    .RESET_B(_0469_),
    .Q(\output_c[12][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5234_ (.CLK(clknet_leaf_10_clk),
    .D(_0999_),
    .RESET_B(_0470_),
    .Q(\output_c[12][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5235_ (.CLK(clknet_leaf_10_clk),
    .D(_1000_),
    .RESET_B(_0471_),
    .Q(\output_c[12][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5236_ (.CLK(clknet_leaf_8_clk),
    .D(_1001_),
    .RESET_B(_0472_),
    .Q(\output_c[12][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5237_ (.CLK(clknet_leaf_14_clk),
    .D(_1002_),
    .RESET_B(_0473_),
    .Q(\output_c[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5238_ (.CLK(clknet_leaf_5_clk),
    .D(_1003_),
    .RESET_B(_0474_),
    .Q(\output_c[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5239_ (.CLK(clknet_leaf_5_clk),
    .D(_1004_),
    .RESET_B(_0475_),
    .Q(\output_c[13][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5240_ (.CLK(clknet_leaf_5_clk),
    .D(_1005_),
    .RESET_B(_0476_),
    .Q(\output_c[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5241_ (.CLK(clknet_leaf_6_clk),
    .D(_1006_),
    .RESET_B(_0477_),
    .Q(\output_c[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5242_ (.CLK(clknet_leaf_6_clk),
    .D(_1007_),
    .RESET_B(_0478_),
    .Q(\output_c[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5243_ (.CLK(clknet_leaf_6_clk),
    .D(_1008_),
    .RESET_B(_0479_),
    .Q(\output_c[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5244_ (.CLK(clknet_leaf_6_clk),
    .D(_1009_),
    .RESET_B(_0480_),
    .Q(\output_c[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5245_ (.CLK(clknet_leaf_7_clk),
    .D(_1010_),
    .RESET_B(_0481_),
    .Q(\output_c[13][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5246_ (.CLK(clknet_leaf_7_clk),
    .D(_1011_),
    .RESET_B(_0482_),
    .Q(\output_c[13][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5247_ (.CLK(clknet_leaf_7_clk),
    .D(_1012_),
    .RESET_B(_0483_),
    .Q(\output_c[13][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5248_ (.CLK(clknet_leaf_1_clk),
    .D(_1013_),
    .RESET_B(_0484_),
    .Q(\output_c[13][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5249_ (.CLK(clknet_leaf_1_clk),
    .D(_1014_),
    .RESET_B(_0485_),
    .Q(\output_c[13][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5250_ (.CLK(clknet_leaf_1_clk),
    .D(_1015_),
    .RESET_B(_0486_),
    .Q(\output_c[13][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5251_ (.CLK(clknet_leaf_1_clk),
    .D(_1016_),
    .RESET_B(_0487_),
    .Q(\output_c[13][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5252_ (.CLK(clknet_leaf_1_clk),
    .D(_1017_),
    .RESET_B(_0488_),
    .Q(\output_c[13][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5253_ (.CLK(clknet_leaf_1_clk),
    .D(_1018_),
    .RESET_B(_0489_),
    .Q(\output_c[13][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5254_ (.CLK(clknet_leaf_1_clk),
    .D(_1019_),
    .RESET_B(_0490_),
    .Q(\output_c[13][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5255_ (.CLK(clknet_leaf_1_clk),
    .D(_1020_),
    .RESET_B(_0491_),
    .Q(\output_c[13][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5256_ (.CLK(clknet_leaf_1_clk),
    .D(_1021_),
    .RESET_B(_0492_),
    .Q(\output_c[13][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5257_ (.CLK(clknet_leaf_0_clk),
    .D(_1022_),
    .RESET_B(_0493_),
    .Q(\output_c[13][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5258_ (.CLK(clknet_leaf_1_clk),
    .D(_1023_),
    .RESET_B(_0494_),
    .Q(\output_c[13][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5259_ (.CLK(clknet_leaf_0_clk),
    .D(_1024_),
    .RESET_B(_0495_),
    .Q(\output_c[13][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5260_ (.CLK(clknet_leaf_0_clk),
    .D(_1025_),
    .RESET_B(_0496_),
    .Q(\output_c[13][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5261_ (.CLK(clknet_leaf_2_clk),
    .D(_1026_),
    .RESET_B(_0497_),
    .Q(\output_c[13][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5262_ (.CLK(clknet_leaf_2_clk),
    .D(_1027_),
    .RESET_B(_0498_),
    .Q(\output_c[13][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5263_ (.CLK(clknet_leaf_1_clk),
    .D(_1028_),
    .RESET_B(_0499_),
    .Q(\output_c[13][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5264_ (.CLK(clknet_leaf_1_clk),
    .D(_1029_),
    .RESET_B(_0500_),
    .Q(\output_c[13][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5265_ (.CLK(clknet_leaf_1_clk),
    .D(_1030_),
    .RESET_B(_0501_),
    .Q(\output_c[13][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5266_ (.CLK(clknet_leaf_1_clk),
    .D(_1031_),
    .RESET_B(_0502_),
    .Q(\output_c[13][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5267_ (.CLK(clknet_leaf_2_clk),
    .D(_1032_),
    .RESET_B(_0503_),
    .Q(\output_c[13][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5268_ (.CLK(clknet_leaf_2_clk),
    .D(_1033_),
    .RESET_B(_0504_),
    .Q(\output_c[13][31] ));
 sky130_fd_sc_hd__dfrtp_1 _5269_ (.CLK(clknet_leaf_4_clk),
    .D(_1034_),
    .RESET_B(_0505_),
    .Q(\output_c[14][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5270_ (.CLK(clknet_leaf_4_clk),
    .D(_1035_),
    .RESET_B(_0506_),
    .Q(\output_c[14][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5271_ (.CLK(clknet_leaf_3_clk),
    .D(_1036_),
    .RESET_B(_0507_),
    .Q(\output_c[14][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5272_ (.CLK(clknet_leaf_3_clk),
    .D(_1037_),
    .RESET_B(_0508_),
    .Q(\output_c[14][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5273_ (.CLK(clknet_leaf_2_clk),
    .D(_1038_),
    .RESET_B(_0509_),
    .Q(\output_c[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5274_ (.CLK(clknet_leaf_2_clk),
    .D(_1039_),
    .RESET_B(_0510_),
    .Q(\output_c[14][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5275_ (.CLK(clknet_leaf_2_clk),
    .D(_1040_),
    .RESET_B(_0511_),
    .Q(\output_c[14][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5276_ (.CLK(clknet_leaf_2_clk),
    .D(_1041_),
    .RESET_B(_0512_),
    .Q(\output_c[14][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5277_ (.CLK(clknet_leaf_2_clk),
    .D(_1042_),
    .RESET_B(_0513_),
    .Q(\output_c[14][8] ));
 sky130_fd_sc_hd__dfrtp_1 _5278_ (.CLK(clknet_leaf_2_clk),
    .D(_1043_),
    .RESET_B(_0514_),
    .Q(\output_c[14][9] ));
 sky130_fd_sc_hd__dfrtp_1 _5279_ (.CLK(clknet_leaf_2_clk),
    .D(_1044_),
    .RESET_B(_0515_),
    .Q(\output_c[14][10] ));
 sky130_fd_sc_hd__dfrtp_1 _5280_ (.CLK(clknet_leaf_2_clk),
    .D(_1045_),
    .RESET_B(_0516_),
    .Q(\output_c[14][11] ));
 sky130_fd_sc_hd__dfrtp_1 _5281_ (.CLK(clknet_leaf_3_clk),
    .D(_1046_),
    .RESET_B(_0517_),
    .Q(\output_c[14][12] ));
 sky130_fd_sc_hd__dfrtp_1 _5282_ (.CLK(clknet_leaf_0_clk),
    .D(_1047_),
    .RESET_B(_0518_),
    .Q(\output_c[14][13] ));
 sky130_fd_sc_hd__dfrtp_1 _5283_ (.CLK(clknet_leaf_0_clk),
    .D(_1048_),
    .RESET_B(_0519_),
    .Q(\output_c[14][14] ));
 sky130_fd_sc_hd__dfrtp_1 _5284_ (.CLK(clknet_leaf_37_clk),
    .D(_1049_),
    .RESET_B(_0520_),
    .Q(\output_c[14][15] ));
 sky130_fd_sc_hd__dfrtp_1 _5285_ (.CLK(clknet_leaf_3_clk),
    .D(_1050_),
    .RESET_B(_0521_),
    .Q(\output_c[14][16] ));
 sky130_fd_sc_hd__dfrtp_1 _5286_ (.CLK(clknet_leaf_37_clk),
    .D(_1051_),
    .RESET_B(_0522_),
    .Q(\output_c[14][17] ));
 sky130_fd_sc_hd__dfrtp_1 _5287_ (.CLK(clknet_leaf_37_clk),
    .D(_1052_),
    .RESET_B(_0523_),
    .Q(\output_c[14][18] ));
 sky130_fd_sc_hd__dfrtp_1 _5288_ (.CLK(clknet_leaf_37_clk),
    .D(_1053_),
    .RESET_B(_0524_),
    .Q(\output_c[14][19] ));
 sky130_fd_sc_hd__dfrtp_1 _5289_ (.CLK(clknet_leaf_3_clk),
    .D(_1054_),
    .RESET_B(_0525_),
    .Q(\output_c[14][20] ));
 sky130_fd_sc_hd__dfrtp_1 _5290_ (.CLK(clknet_leaf_36_clk),
    .D(_1055_),
    .RESET_B(_0526_),
    .Q(\output_c[14][21] ));
 sky130_fd_sc_hd__dfrtp_1 _5291_ (.CLK(clknet_leaf_36_clk),
    .D(_1056_),
    .RESET_B(_0527_),
    .Q(\output_c[14][22] ));
 sky130_fd_sc_hd__dfrtp_1 _5292_ (.CLK(clknet_leaf_4_clk),
    .D(_1057_),
    .RESET_B(_0528_),
    .Q(\output_c[14][23] ));
 sky130_fd_sc_hd__dfrtp_1 _5293_ (.CLK(clknet_leaf_3_clk),
    .D(_1058_),
    .RESET_B(_0529_),
    .Q(\output_c[14][24] ));
 sky130_fd_sc_hd__dfrtp_1 _5294_ (.CLK(clknet_leaf_4_clk),
    .D(_1059_),
    .RESET_B(_0530_),
    .Q(\output_c[14][25] ));
 sky130_fd_sc_hd__dfrtp_1 _5295_ (.CLK(clknet_leaf_4_clk),
    .D(_1060_),
    .RESET_B(_0531_),
    .Q(\output_c[14][26] ));
 sky130_fd_sc_hd__dfrtp_1 _5296_ (.CLK(clknet_leaf_2_clk),
    .D(_1061_),
    .RESET_B(_0532_),
    .Q(\output_c[14][27] ));
 sky130_fd_sc_hd__dfrtp_1 _5297_ (.CLK(clknet_leaf_2_clk),
    .D(_1062_),
    .RESET_B(_0533_),
    .Q(\output_c[14][28] ));
 sky130_fd_sc_hd__dfrtp_1 _5298_ (.CLK(clknet_leaf_6_clk),
    .D(_1063_),
    .RESET_B(_0534_),
    .Q(\output_c[14][29] ));
 sky130_fd_sc_hd__dfrtp_1 _5299_ (.CLK(clknet_leaf_6_clk),
    .D(_1064_),
    .RESET_B(_0535_),
    .Q(\output_c[14][30] ));
 sky130_fd_sc_hd__dfrtp_1 _5300_ (.CLK(clknet_leaf_6_clk),
    .D(_1065_),
    .RESET_B(_0536_),
    .Q(\output_c[14][31] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_785 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(input_a_serial),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(rst),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 output3 (.A(net3),
    .X(output_c_serial[0]));
 sky130_fd_sc_hd__clkbuf_4 output4 (.A(net4),
    .X(output_c_serial[10]));
 sky130_fd_sc_hd__clkbuf_4 output5 (.A(net5),
    .X(output_c_serial[11]));
 sky130_fd_sc_hd__clkbuf_4 output6 (.A(net6),
    .X(output_c_serial[12]));
 sky130_fd_sc_hd__clkbuf_4 output7 (.A(net7),
    .X(output_c_serial[13]));
 sky130_fd_sc_hd__clkbuf_4 output8 (.A(net8),
    .X(output_c_serial[14]));
 sky130_fd_sc_hd__clkbuf_4 output9 (.A(net9),
    .X(output_c_serial[15]));
 sky130_fd_sc_hd__clkbuf_4 output10 (.A(net10),
    .X(output_c_serial[16]));
 sky130_fd_sc_hd__clkbuf_4 output11 (.A(net11),
    .X(output_c_serial[17]));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(output_c_serial[18]));
 sky130_fd_sc_hd__clkbuf_4 output13 (.A(net13),
    .X(output_c_serial[19]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(output_c_serial[1]));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(output_c_serial[20]));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(output_c_serial[21]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(output_c_serial[22]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(output_c_serial[23]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(output_c_serial[24]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(output_c_serial[25]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(output_c_serial[26]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(output_c_serial[27]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(output_c_serial[28]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(output_c_serial[29]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(output_c_serial[2]));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net26),
    .X(output_c_serial[30]));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net27),
    .X(output_c_serial[31]));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net28),
    .X(output_c_serial[3]));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net29),
    .X(output_c_serial[4]));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net30),
    .X(output_c_serial[5]));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net31),
    .X(output_c_serial[6]));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net32),
    .X(output_c_serial[7]));
 sky130_fd_sc_hd__clkbuf_4 output33 (.A(net33),
    .X(output_c_serial[8]));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net34),
    .X(output_c_serial[9]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\output_c[6][31] ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\output_c[1][31] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\output_c[10][31] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\output_c[4][31] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\output_c[11][31] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\output_c[8][31] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\output_c[12][31] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\output_c[2][31] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\output_c[9][31] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\output_c[13][31] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\output_c[3][31] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0713_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\output_c[5][31] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\output_c[0][31] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\output_c[7][31] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\output_c[15][31] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\output_c[10][15] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\output_c[3][15] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\output_c[12][15] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\output_c[9][15] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\output_c[6][15] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\output_c[8][15] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\output_c[2][15] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\output_c[14][31] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\output_c[1][30] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\state[0] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\output_c[5][15] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\output_c[12][30] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\output_c[13][15] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\output_c[15][15] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\output_c[4][15] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\output_c[0][15] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\output_c[15][23] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\output_c[7][15] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\output_c[7][25] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\output_c[10][30] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\output_c[11][15] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\output_c[11][30] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\output_c[13][30] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\output_c[1][25] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\output_c[6][30] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\output_c[9][30] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\output_c[15][30] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\output_c[8][25] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\output_c[1][15] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\output_c[2][30] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\output_c[4][30] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\output_c[8][30] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\output_c[7][30] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\output_c[5][30] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\output_c[3][30] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0712_),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\output_c[12][19] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\output_c[14][24] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\output_c[11][23] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\output_c[0][30] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\output_c[14][7] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\output_c[3][10] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\output_c[14][23] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\output_c[9][11] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_1466_),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\output_c[0][22] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\output_c[11][26] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\output_c[13][11] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_1208_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\output_c[3][22] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\output_c[1][22] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\output_c[6][11] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_1650_),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\output_c[14][27] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\output_c[8][10] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\output_c[4][10] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\output_c[7][11] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_1587_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\output_c[10][26] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\output_c[9][22] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\output_c[4][11] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\output_c[11][11] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_1335_),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\output_c[4][20] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\output_c[15][11] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_2137_),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\output_c[1][27] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_1938_),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\output_c[2][10] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\output_c[4][26] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\output_c[5][10] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\output_c[15][10] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\output_c[6][19] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\output_c[2][11] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\output_c[6][22] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\output_c[11][27] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\output_c[0][10] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\output_c[9][10] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\output_c[14][19] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\output_c[12][20] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\output_c[4][21] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\output_c[11][18] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\output_c[5][11] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\output_c[3][19] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\output_c[13][19] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\output_c[15][18] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\output_c[9][26] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\output_c[12][10] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\output_c[6][10] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\output_c[7][26] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\output_c[8][11] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\output_c[11][0] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\output_c[12][11] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\output_c[15][22] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0560_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\output_c[0][11] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\output_c[9][19] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\output_c[7][18] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\output_c[12][23] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_1253_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\output_c[7][22] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\output_c[5][22] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\output_c[14][15] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\output_c[11][20] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\output_c[9][0] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\output_c[10][11] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_1401_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\output_c[0][18] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\output_c[11][10] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\output_c[2][22] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\output_c[7][10] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\output_c[1][26] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\output_c[13][23] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_1190_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\output_c[2][3] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\output_c[13][26] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\output_c[1][0] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\output_c[10][0] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\output_c[1][3] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\output_c[3][6] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\output_c[1][18] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\output_c[12][22] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\output_c[12][0] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\output_c[10][10] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\output_c[15][26] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\output_c[13][22] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\output_c[0][0] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\output_c[13][10] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\output_c[3][11] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\output_c[5][0] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\output_c[10][22] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\output_c[10][18] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\output_c[3][0] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\output_c[2][0] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\output_c[8][16] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\output_c[12][26] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\output_c[5][9] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_1715_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\output_c[2][19] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\output_c[4][18] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\output_c[6][0] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\output_c[14][30] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_1087_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\output_c[13][0] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\output_c[3][21] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_1820_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\output_c[9][3] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0877_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\output_c[8][18] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\output_c[0][3] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\output_c[12][13] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\output_c[8][27] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_1504_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\output_c[10][9] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_1402_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\output_c[10][14] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\output_c[4][1] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\output_c[8][0] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\output_c[3][26] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\output_c[10][16] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\output_c[7][27] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\output_c[1][10] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\output_c[6][26] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\output_c[12][18] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_1260_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\output_c[7][0] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\output_c[1][16] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\output_c[8][3] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\output_c[1][11] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\output_c[8][22] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\output_c[1][21] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_1947_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\output_c[5][19] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\output_c[5][14] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\output_c[15][0] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\output_c[3][3] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\output_c[11][3] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\output_c[6][18] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_1638_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\output_c[9][13] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\output_c[5][26] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\output_c[11][13] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\output_c[4][0] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\output_c[10][20] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\output_c[3][14] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\output_c[13][20] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\output_c[0][16] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\output_c[9][14] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\output_c[6][8] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\output_c[4][13] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\output_c[7][16] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\output_c[3][16] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\output_c[6][21] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_1635_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\output_c[3][13] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\output_c[9][17] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\output_c[10][21] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\output_c[2][26] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\output_c[7][3] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\output_c[5][8] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\output_c[3][8] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\output_c[10][8] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\output_c[8][9] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_1528_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\output_c[15][3] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\output_c[3][28] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\output_c[15][27] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\output_c[3][20] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\output_c[8][26] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\output_c[10][28] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\output_c[3][9] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\output_c[1][6] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\output_c[3][29] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\output_c[12][3] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\output_c[9][28] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\output_c[1][20] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\output_c[14][29] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\output_c[13][6] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\output_c[12][17] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\output_c[8][8] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\output_c[7][13] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\output_c[15][8] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\output_c[8][28] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\output_c[6][6] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\output_c[13][28] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\output_c[9][6] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\output_c[2][14] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\output_c[3][17] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\output_c[13][13] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\output_c[9][20] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\output_c[7][9] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_1588_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\output_c[12][1] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\output_c[2][21] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_1883_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\output_c[6][3] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\output_c[8][6] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\output_c[11][14] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\output_c[4][3] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\output_c[9][9] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_1467_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\output_c[7][12] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\output_c[11][22] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\output_c[13][14] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\output_c[10][12] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\output_c[12][28] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\output_c[13][17] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\output_c[0][8] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\output_c[6][20] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\output_c[7][6] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\output_c[6][17] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\output_c[4][9] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_1776_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\output_c[14][22] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\output_c[9][8] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\output_c[9][18] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\output_c[15][25] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\output_c[12][8] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\output_c[12][6] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\output_c[2][13] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\output_c[15][13] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\output_c[5][28] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\output_c[12][9] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\output_c[5][20] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\output_c[4][8] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\output_c[5][29] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_0775_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\output_c[9][29] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0903_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\output_c[15][1] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\output_c[10][29] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\output_c[3][18] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\output_c[6][13] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\output_c[4][6] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\output_c[9][12] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\output_c[12][16] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\output_c[0][20] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\output_c[11][8] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\output_c[0][26] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\output_c[9][1] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\output_c[2][20] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\output_c[0][13] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\output_c[8][29] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\output_c[13][18] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\output_c[11][6] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\output_c[11][28] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\output_c[7][20] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\output_c[15][28] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\output_c[13][8] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\output_c[5][13] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\output_c[2][12] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\output_c[1][29] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_1934_),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\output_c[15][14] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\output_c[2][28] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\output_c[9][21] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\output_c[2][8] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\output_c[5][1] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\output_c[11][24] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\output_c[2][2] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0652_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\output_c[7][21] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\output_c[14][11] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\output_c[10][13] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\output_c[6][9] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\output_c[2][17] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\output_c[2][6] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\output_c[10][6] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\output_c[1][28] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\output_c[8][12] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\output_c[0][21] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\output_c[4][29] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_1747_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\output_c[7][8] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\output_c[5][6] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\output_c[4][22] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\output_c[6][1] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\output_c[4][28] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\output_c[12][12] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\output_c[11][25] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\output_c[5][3] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\output_c[2][18] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\output_c[4][14] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\output_c[11][17] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\output_c[1][1] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\output_c[2][9] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\output_c[2][1] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\output_c[1][8] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\output_c[0][6] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\output_c[12][29] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\output_c[11][1] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\output_c[15][17] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\output_c[13][9] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\output_c[8][1] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\output_c[11][29] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\output_c[5][17] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\output_c[6][29] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_1620_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\output_c[3][12] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\output_c[0][28] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\output_c[13][12] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\output_c[6][12] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\output_c[0][1] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\output_c[13][29] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\output_c[13][3] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\output_c[13][1] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\output_c[4][17] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\output_c[6][14] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\output_c[7][28] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\output_c[15][29] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\output_c[11][16] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\output_c[4][23] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\output_c[1][9] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\output_c[10][3] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\output_c[15][9] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\output_c[7][1] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\output_c[1][13] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\output_c[12][2] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\output_c[0][14] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\output_c[3][1] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\output_c[11][9] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\output_c[6][28] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\output_c[0][2] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0588_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\output_c[8][20] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\output_c[0][9] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\output_c[5][21] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\output_c[13][2] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\output_c[14][12] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\output_c[15][12] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\output_c[15][2] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\output_c[0][12] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\output_c[5][18] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\output_c[11][2] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0940_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\output_c[15][20] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\output_c[15][6] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\output_c[8][2] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_0844_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\output_c[2][29] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\output_c[8][13] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\output_c[7][29] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\output_c[1][12] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\output_c[14][16] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\output_c[0][29] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\output_c[10][1] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\output_c[8][21] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\output_c[4][2] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_0716_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\output_c[5][2] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\output_c[11][12] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\output_c[1][2] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_0620_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\output_c[4][16] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\output_c[3][2] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\output_c[9][2] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(_0876_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\output_c[13][16] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\output_c[12][5] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\output_c[6][2] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_0780_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\output_c[14][1] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\output_c[7][5] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\output_c[14][14] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\output_c[9][5] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\output_c[6][5] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\output_c[4][12] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\output_c[12][14] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\output_c[5][12] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\output_c[11][5] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\output_c[13][5] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\output_c[10][2] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\output_c[2][5] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\output_c[14][6] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\output_c[14][8] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\output_c[8][5] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\output_c[14][3] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\output_c[4][5] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\output_c[8][17] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\output_c[15][5] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\output_c[5][5] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\output_c[7][2] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\output_c[0][5] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\output_c[4][25] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\output_c[1][5] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\output_c[10][17] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\output_c[14][18] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\output_c[14][26] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\output_c[0][17] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\output_c[10][5] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\output_c[1][17] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\output_c[3][5] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\output_c[7][17] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\output_c[8][23] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\output_c[10][23] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\output_c[1][23] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_1944_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\output_c[7][23] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\output_c[0][23] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\input_a[15] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\output_c[5][28] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\output_c[11][25] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\output_c[10][30] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\output_c[15][25] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\output_c[12][30] ),
    .X(net495));
endmodule
