VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO matrix_mult3
  CLASS BLOCK ;
  FOREIGN matrix_mult3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 220.665 BY 231.385 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 220.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 220.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 215.060 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 215.060 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 220.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 220.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 215.060 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 215.060 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END clk
  PIN input_a_serial
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 227.385 113.070 231.385 ;
    END
  END input_a_serial
  PIN input_b_serial
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END input_b_serial
  PIN output_c_serial[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END output_c_serial[0]
  PIN output_c_serial[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END output_c_serial[10]
  PIN output_c_serial[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END output_c_serial[11]
  PIN output_c_serial[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END output_c_serial[12]
  PIN output_c_serial[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END output_c_serial[13]
  PIN output_c_serial[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END output_c_serial[14]
  PIN output_c_serial[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END output_c_serial[15]
  PIN output_c_serial[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END output_c_serial[16]
  PIN output_c_serial[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END output_c_serial[17]
  PIN output_c_serial[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END output_c_serial[18]
  PIN output_c_serial[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END output_c_serial[19]
  PIN output_c_serial[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END output_c_serial[1]
  PIN output_c_serial[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END output_c_serial[20]
  PIN output_c_serial[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END output_c_serial[21]
  PIN output_c_serial[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END output_c_serial[22]
  PIN output_c_serial[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END output_c_serial[23]
  PIN output_c_serial[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END output_c_serial[24]
  PIN output_c_serial[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END output_c_serial[25]
  PIN output_c_serial[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END output_c_serial[26]
  PIN output_c_serial[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END output_c_serial[27]
  PIN output_c_serial[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END output_c_serial[28]
  PIN output_c_serial[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END output_c_serial[29]
  PIN output_c_serial[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END output_c_serial[2]
  PIN output_c_serial[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END output_c_serial[30]
  PIN output_c_serial[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END output_c_serial[31]
  PIN output_c_serial[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END output_c_serial[3]
  PIN output_c_serial[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END output_c_serial[4]
  PIN output_c_serial[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END output_c_serial[5]
  PIN output_c_serial[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END output_c_serial[6]
  PIN output_c_serial[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END output_c_serial[7]
  PIN output_c_serial[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END output_c_serial[8]
  PIN output_c_serial[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END output_c_serial[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END rst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 214.820 220.405 ;
      LAYER met1 ;
        RECT 4.670 9.900 215.120 220.560 ;
      LAYER met2 ;
        RECT 4.690 227.105 112.510 227.385 ;
        RECT 113.350 227.105 213.340 227.385 ;
        RECT 4.690 4.280 213.340 227.105 ;
        RECT 4.690 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 86.750 4.280 ;
        RECT 87.590 4.000 89.970 4.280 ;
        RECT 90.810 4.000 93.190 4.280 ;
        RECT 94.030 4.000 96.410 4.280 ;
        RECT 97.250 4.000 213.340 4.280 ;
      LAYER met3 ;
        RECT 3.990 215.240 211.535 220.485 ;
        RECT 4.400 213.840 211.535 215.240 ;
        RECT 3.990 140.440 211.535 213.840 ;
        RECT 4.400 139.040 211.535 140.440 ;
        RECT 3.990 137.040 211.535 139.040 ;
        RECT 4.400 135.640 211.535 137.040 ;
        RECT 3.990 133.640 211.535 135.640 ;
        RECT 4.400 132.240 211.535 133.640 ;
        RECT 3.990 130.240 211.535 132.240 ;
        RECT 4.400 128.840 211.535 130.240 ;
        RECT 3.990 126.840 211.535 128.840 ;
        RECT 4.400 125.440 211.535 126.840 ;
        RECT 3.990 123.440 211.535 125.440 ;
        RECT 4.400 122.040 211.535 123.440 ;
        RECT 3.990 120.040 211.535 122.040 ;
        RECT 4.400 118.640 211.535 120.040 ;
        RECT 3.990 116.640 211.535 118.640 ;
        RECT 4.400 115.240 211.535 116.640 ;
        RECT 3.990 113.240 211.535 115.240 ;
        RECT 4.400 111.840 211.535 113.240 ;
        RECT 3.990 109.840 211.535 111.840 ;
        RECT 4.400 108.440 211.535 109.840 ;
        RECT 3.990 106.440 211.535 108.440 ;
        RECT 4.400 105.040 211.535 106.440 ;
        RECT 3.990 103.040 211.535 105.040 ;
        RECT 4.400 101.640 211.535 103.040 ;
        RECT 3.990 99.640 211.535 101.640 ;
        RECT 4.400 98.240 211.535 99.640 ;
        RECT 3.990 96.240 211.535 98.240 ;
        RECT 4.400 94.840 211.535 96.240 ;
        RECT 3.990 92.840 211.535 94.840 ;
        RECT 4.400 91.440 211.535 92.840 ;
        RECT 3.990 89.440 211.535 91.440 ;
        RECT 4.400 88.040 211.535 89.440 ;
        RECT 3.990 86.040 211.535 88.040 ;
        RECT 4.400 84.640 211.535 86.040 ;
        RECT 3.990 82.640 211.535 84.640 ;
        RECT 4.400 81.240 211.535 82.640 ;
        RECT 3.990 79.240 211.535 81.240 ;
        RECT 4.400 77.840 211.535 79.240 ;
        RECT 3.990 75.840 211.535 77.840 ;
        RECT 4.400 74.440 211.535 75.840 ;
        RECT 3.990 72.440 211.535 74.440 ;
        RECT 4.400 71.040 211.535 72.440 ;
        RECT 3.990 69.040 211.535 71.040 ;
        RECT 4.400 67.640 211.535 69.040 ;
        RECT 3.990 65.640 211.535 67.640 ;
        RECT 4.400 64.240 211.535 65.640 ;
        RECT 3.990 62.240 211.535 64.240 ;
        RECT 4.400 60.840 211.535 62.240 ;
        RECT 3.990 10.715 211.535 60.840 ;
      LAYER met4 ;
        RECT 26.975 13.095 174.240 131.745 ;
        RECT 176.640 13.095 177.540 131.745 ;
        RECT 179.940 13.095 193.825 131.745 ;
  END
END matrix_mult3
END LIBRARY

